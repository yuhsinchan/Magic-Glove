`include "Top.sv"
//`include "Random.sv"
`include "DE2_115/PreviousValue.sv"
`include "DE2_115/SevenHexDecoder.sv"
`include "DE2_115/Debounce.sv"
`include "DE2_115/DE2_115.sv"

`timescale 1ns / 100ps
module Dictionary(
	input          i_clk,
	input          i_rst_n,
	input          i_start,
	input  [119:0] i_word,
	output         o_finish,
	output [119:0] o_word,
	output [1:0]   o_state,
	output [119:0] o_DTW_candidate_word [0:19]
);
	parameter DICT_SIZE = 500;
	localparam bit [119:0] dict [0:DICT_SIZE - 1] = '{
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100100000111100010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000100000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000111000000001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000111100000110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000010000100000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011000010010000100000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000101000000100100010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000111100011001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000111100001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010001001000000001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000011110001001000000110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000101010000111100011001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000110000000001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000101100000000100001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110000010100001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000100100000111100001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110000000100010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011000000100100010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000011010000111100001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010101000011110000001000000001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001110000000100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110000000100001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000001100010010000000010000010100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001010001001000000110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001010100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100001010100001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000111000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000101000010000001010000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100001110,
		120'b000000000000000000000000000000000000111000001111000010010001010000000001000011010001001000001111000001100000111000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000011010000100100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000001010000100000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000101000000100100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010000000100001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000010000100000010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000011000010010000100000010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000001001000001010000100000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011000101110000010100001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001010100001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010001001100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010000111000000001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010010000001010000100000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000011000000111000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110000100100001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000001010000100000010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000010100000000110000000100010100000011100000111100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000100100000010100001000,
		120'b000000000000000000000000000000000000000000000000000000000001001100010011000001010000111000001001000100110001010100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000100000010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010100010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000100110000110000000001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110000111100001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000011000000010100001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000010100000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111000001010000100100010110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010000111000001001000011000000111000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010011000100100000100100000110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100000001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000001010000010100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001100000101010000111100010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110000111100001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000100100000010100010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011,
		120'b000000000000000000000000000000000000000000000000000000000001001100000101000000110000100100010110000100100000010100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000011010000111100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010011000001010000100000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100000011000010010000110000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110001010000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000010110000100100001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000101000000110000100100010110000100100000010100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000010000100000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011100000100100000110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000011000010010001001000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000101000000000100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000000110000000100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000111100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010000110000010000000011110000010100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100110000100100001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000011010000000100001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100110001010100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000001010001011000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010100000000010001010000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000010000010100011001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010000000100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000101000000111000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001001000000010000110100000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110001011100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000001010000001100000000010000010100001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001100000100100000111100010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000110000000010100001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001010001001100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000100100000111100010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100110000000100001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100110000111100001101,
		120'b000000000000000000000000000000000000000000000000000000000001001100010100000000110001010100000100000011110001001000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100001001000100110001010100001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010001010100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000101000000000100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000010110000000100001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000001010000100000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000110000010101000011110000100000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000010100000000110001010100000100000011110001001000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000011010000010100010100000100110001100100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100110000111100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000010100001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000101000000100100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000110010000001100001001000011000000111100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000100100000010100000010000011010001010100001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000110001010100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010001001100000001000001010000110000010000,
		120'b000000000000000000000000000000000000000000000000000001010000110000000010000000010000110000001001000000010001011000000001,
		120'b000000000000000000000000000000000000000000000000000101000000100000000111000010010001001000011001000100000000111100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000010100000100100000111100010000000100000001010100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000101000001110000000100010011000100110000010100001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000101000101000000011000000001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100110000010100000010,
		120'b000000000000000000000000000000000000000000000000000000000000010100010010000000010001011100010100000001100000111100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000001010000100000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011110000111100000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000101000001000000100100010110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011000000010100010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010010000001010000100000010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000001100000111000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110001010000001000000001110000100100010010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000110000100100001100000000100001010100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100001011000011110000111100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001110000100100001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000011000000111100001111000010000000001100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000001000000001110001010100001111000100100000100000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000110000000100000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100001011000011100000100100001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000100000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000101110000010100001001000101100000010100010010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100010010000000010000010100011001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000101000001000001001000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000100100000010100010110,
		120'b000000000000000000000000000000000000000000000000000000000000000000011001000000110000000100010110000010010001001000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000011110000111100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100001101000001010001010000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000011001000011100000000100010000000011010000111100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000010100010010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010101000011110001001000000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000010100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001010000010100001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000011100000000100001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000001010001001100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010010000000100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011000001010000111100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000010100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000101000001000000111000010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000001100000000010001001000000101000011100000010100000111,
		120'b000000000000000000000000000000000000000000000000000000000000100000000011000100100000000100000101000100110000010100010010,
		120'b000000000000000000000000000000000000000000011001000101000000100100010011000100100000010100010110000010010000111000010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000011001000100100000000100010101000011100000000100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000010010000000100001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011000001010100000110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000010011000101110000010100001001000101100000010100010010,
		120'b000000000000000000000000000000000000000000000000000000000000000000001101000000010001001000000111000011110001001000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001100000100100001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111000011110000111000001011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000101000011010000000100000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010000000100010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011000110010000000100000100,
		120'b000000000000000000000000000000000000000000010100000011100000010100001101000001010000011100000001000011100000000100001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100100000000100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001100000101010000111100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000001000001010001001000000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000010100010100000010010000111000010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000101000101000000111100001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000010000010100010010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000001010001010000001001,
		120'b000000000000000000001100000000010000111000001111000010010001010000000001000011100001001000000101000101000000111000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000100100000010100010100000011100000010100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000000010000001000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100110001010100001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010010000011110001010000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000011000000010100010110000000010001001000010100,
		120'b000000000000000000000000000000000000000000000000000000000001001100010100000011100000010100001101000011010000111100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001000000000100001101,
		120'b000000000000000000000000000000000001010000001110000001010000110100010000000011110000110000000101000101100000010100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000001001000001111000100000000010100010010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000100100000010100000010000011010000010100001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000010011000011000000100100000001000101000000010100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000011100000100100001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100001101000100100000010100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010001001000001111000001100000010100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110000110000000101000101000000111100001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011100000010100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000001000000001110000100100010010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000100000001100100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000101000100110001010100000001000000110000010100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000001000000110000111100001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010011000011110000100000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001110000010010001001100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000010011000101000000110000010101000100110000010100010010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010000001100001001000001100000011000001111,
		120'b000000000000000000000000000000000000000000000000000011100000111100001001000101000000000100000011000101010000010000000101,
		120'b000000000000000000000000000000000000000000000000000000000000110000000001000011100000111100001001000101000000000100001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000011100000011100001001000100110000010100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000010110000000100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000010100010100000100110000111100010000,
		120'b000000000000000000000000000000000000000000000000000000000001010000000101000011100001001000000101000101000000111000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000010011000100110000010100010010000001000000010000000001,
		120'b000000000000000000000000000000000000000000000000000110010001010000001001000011100001010100001101000011010000111100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000011100000100100001000000101000000100100010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110000010100010100000000010001010000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001010001001000000001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000011100000000100010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001110000011110000100000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001011000000100,
		120'b000000000000000000000000000000000000000000000000000000000000011100001110000010010001000000010000000010010000100000010011,
		120'b000000000000000000000000000000000000000000000000000000000000010000000101000101100001001000000101000100110000010100010010,
		120'b000000000000000000000000000000000000000000000000000000000000000000010100000000110000010100001010000000100001010100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000001110000001010000010100010111000101000000010100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100010101000100100000111100000110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000110010000110000001001000011010000000100000110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011100000111100001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000101000100110000000100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001000000111100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111000011110000100000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000001010001011000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100000011000000010000110000000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100000011000001010000100000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000001100000000010000100100000011000001010001000000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110000010100000011000010010001001000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000101000101000000100100010011000000100000010100010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000101000001000000111000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001110000010010000010100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000101000011010000111100010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000110001010100001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000001110000100100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000011000000100100000110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000011100000100100001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000001010001000000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100000001000001000000111100010100,
		120'b000000000000000000000000000000000000000000011001000001110000111100001100000011110000111000001000000000110000010100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010100000101010000111100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000100110000000100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000010100000000110000010100001010000011110001001000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000011010000000100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000101000001110000000100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000001110000011110000100100010011000100100000010100010110,
		120'b000000000000000000000000000000000000000000000000000000000000000000001110000011110000100100010100000000110000010100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001011100001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001110000101010000111100000110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110001010000010010000011110001000000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010011000101010000111100001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000100000001010001010000000001000011000000010100010010,
		120'b000000000000000000000000000000000000000000000000000000000001100100010100000010010001001000010101000000110000010100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000101000000111100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000110010001010000001110000101010000111100000011,
		120'b000000000000000000000000000000000000000000000000000000000000111000000001000000110000100100010010000001010000110100000001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100010100000011110000100000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000011010000000100000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000010011000100100000010100000010000011010000010100001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000101000101110000111100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001100000010010000100000010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000100100000000100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000001011000100100000111100010111000101000000010100001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000101110000111100000100,
		120'b000000000000000000000000000000000000000000000000000000000001001000000101000101000001010100010000000011010000111100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000010011000011010000010100010100000100110001100100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000101000100100000100000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000001000101000000111100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000011000000010000110000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000111000000101,
		120'b000000000000000000000000000000000000000000000000000001110000111000001001000101110000111100001100000011000000111100000110,
		120'b000000000000000000000000000000000000000000000000000000000000010000000001000011110000110000001110000101110000111100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010000100100001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000010100000101010000111100001000000101000000100100010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000010100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110001001100000101000000110000001100000001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100001110000010010000100000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010100000100100000111100001110,
		120'b000000000000000000000000000000000000000000000000000100110000010100000011000100100001010100001111000100110000010100010010,
		120'b000000000000000000000000000000000000000000000000000000000000000000010100000011100000010100010010000100100001010100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100010100000100110000111100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000100100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001001000001000000010100001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110000000100001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000001100000011110001001000010100000011100000111100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000101000101000000000100010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000011001000100100000111100010100000100110000100100001000,
		120'b000000000000000000000000000000000000000000000000000000000001001100000101000100100001010100010100000000110000100100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000110100000100100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001001000000001,
		120'b000000000000000000000000000000000000000000000000000000000000110000000001000011100000111100010011000100100000010100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000011000011100000100100010011,
		120'b000000000000000000000000000000000000000000000000000001110000111000001001000001000001010100001100000000110000111000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100000010010001010100000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000011110000100000010011,
		120'b000000000000000000000000000000000000000000000000000110010001001000001111000101000000001100000101000100100000100100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010010000000010000111100000010,
		120'b000000000000000000000000000000000000000000000000000000000000111000001111000010010001010000000001000000110000111100001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010000011100001110000000010000100000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010100000010010000100000010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000110000000010100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001100000000010000110100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001110000111000001001000101000000000100010010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000101000000000100010010,
		120'b000000000000000000000000000000000000000000010100000011100000010100001101000011100001001000000101000101100000111100000111,
		120'b000000000000000000000000000000000000000000000000000000000000111000000101000100100000010000001100000010010000100000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001110000111000001001000100100001010100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001001100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000011100001001000010101000101000000010100010010,
		120'b000000000000000000000000000000000000000000000000000000000001001100010100000011100000010100000100000101010001010000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010110,
		120'b000000000000000000000000000000000000000000000000000000000000011100001110000010010001000000010000000011110000100000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000010100000011100001010100001111000000110000001100000001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000101000011010000100100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000101000101000000100100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000101000101100000010100001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000001100000000010001010000001001000001110000100100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000101000011000000100100000110000011110001001000010000,
		120'b000000000000000000000000000000000000000000000000000000000001001100010101000011110000100100010110000001010001001000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000100100000111100000110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110001010000001110000001010001011000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000101100000111100001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000110000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000010000000111100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000010010000000100001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011000000000100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100010010000101010000111100001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000111000000010000110100001001,
		120'b000000000000000000000000000000000000000000010100000011100000010100001101000101000001001000000001000100000000010100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001100000101000000100100010100,
		120'b000000000000000000000000000000000000111000001111000010010001010000010000000010010001001000000011000100110000010100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000111100001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001,
		120'b000000000000000000000000000000000000000000000000000001010000001100001110000000010001001000010101000100110000111000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000010010000001010000100000010100000011110000111000000001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010000100000010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001100000000010000100000010011,
		120'b000000000000000000000000000000000000000000000000000000000001100100010100000100100000010100010000000011110001001000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100010011000000010000110000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001100000010010001010000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100000101000011100000111100001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000011001000101000000100100001100000000010001010100010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100010010000001010001011000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000111000011100000100100010100000100110000100100001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000010100000011100000010100010100000011100000111100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000011001000100100001010000001110000101010000111100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000101000101000000000100010110000010010001001000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010000110000010100000101000000100100001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000001001000100110000100100010110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000101100000000100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100001100000011110000111100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110000111100001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100001100000100000000010100010010,
		120'b000000000000000000000000000000000000000000000000000000000001001000000101000011010000111100010100000100110001010100000011,
		120'b000000000000000000000000000000000000000000000000000000000001001000000101000000100000110100000101000000110000010100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000101000100100000000100010000000011010000111100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110000010100001001000101100000111100001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000101000001000001010100001100000000110000111000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000101000001110000010100001100000011000000111100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010101000011000000000100010110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000101000011000000001100001001000101000001001000000001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000100100000111100011001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000100001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100100000000100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011000000100000111100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000101000001000000100100010110000011110001001000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011110000111100000110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010000001100010010000101010000111100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000100100000111100001000000101000001010100000001,
		120'b000000000000000000000000000000000000000000000000000101000000111000000101000100100000010100000110000001100000100100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100010011000001010001001000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000010010000000010000010100001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000011000000000100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000111000010101000011110001001000000001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000001110000010010001001000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010001001100010010000101010000111100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000111100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000010000000001000011100000000100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000010011000100110000010100000011000011110001001000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000001010000010100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000011110000111100010010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100000011000011110001010000010011,
		120'b000000000000000000000000000000000000000000000000000000000000011100001110000010010000111000001001000000010001001000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000111100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000000100100000100000001010001001000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000001110000010010000111100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000010010000111100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000101000000110000111000000101000010010000001100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000010100001101,
		120'b000000000000000000000000000000000000000000010011000001010000100100010010000011110000011100000101000101000000000100000011,
		120'b000000000000000000000000000000000000000000000000000000000000010000000101000000110000111000000001000101100000010000000001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100110000010100010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000101000011000000000100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000011110000111100001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000001000000100110000100100001100000001110000111000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000001100000010100001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000000010000010100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010001010000000001000101000001001100000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000111100000010,
		120'b000000000000000000000000000000000000000000010011000011100000111100001001000101000000100100000100000011100000111100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000000001100000101000011000000010100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000010011000101110000111100000100000011100000100100010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110000111100010100000011110000100000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010000000100000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000101000100100000100000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000001010000010100010111,
		120'b000000000000000000000000000000000000000000000000000000000001100100010010000011110000011100000101000101000000000100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000101000000111100001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000101100000100100001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000111000100100000000100001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000011001000100100000010100001100000011000000000100000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001100000000100000000100010100,
		120'b000000000000000000000000000000000000000000000000000000000001001000000101000101000001001100001001000001110000010100010010,
		120'b000000000000000000000000000000000000000000000000000000000000000000010010000001010001011000000101000101110000111100001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000011100001010100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000010010000001010000001000001111000101000000001100001111,
		120'b000000000000000000000000000000000000000000000000000000000001001000000101000000100000110100000101000101100000111100001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000000010100001011000100100000000100001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000011001000100100000000100010010000000100000100100001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000110010000110000001100000000010000010100010010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000011100000111100001001000101000000001100000001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010010000000010001010000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110000010100001001000100100000010100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000101000001000000111100001101,
		120'b000000000000000000000000000000000000000000000000000000000001001100000101000100100001010100010100000000010000010100000110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000100100000001,
		120'b000000000000000000000000000000000000000000000000000000000001100100010010000101000001001100010101000001000000111000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000010000110000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000001000011010001010100001000,
		120'b000000000000000000000000000000000000000000000000000000000000010000000101000001000000100100010110000011110001001000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110000010100011001,
		120'b000000000000000000000000000000000000000000000000000000000000010000000101000100100000100100010101000100010000010100010010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000111000001111000000110000010100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000111100001000,
		120'b000000000000000000000000000000000001001100000101000010010001001000001111000100110001001100000101000000110000001100000001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100110000111100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001001000101100000111100001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110000110100010101000100100000111100000110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000011000100100000000100001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001100,
		120'b000000000000000000000000000000000000000000000000000100100000010100000010000011010000010100010100000100000000010100010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000100100000010100010100000101000000010100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010000000100010011,
		120'b000000000000000000000000000000000000000000000000000100110000111000001111000010010001010000010011000001010001010100010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000011000001010100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100001111000010000000000100011001
	};
	
	localparam S_IDLE = 2'd0;
	localparam S_CALC = 2'd1;
	localparam S_DONE = 2'd2;
	
	logic [1:0] state_r, state_w;
	logic finish_r, finish_w;
	
	logic similarity_start_r, similarity_start_w;
	logic similarity_finish_r, pre_similarity_finish_r;
	logic similarity_finish;
	logic [2:0] DTW_state_r; // debug
	logic DTW_start_r, DTW_start_w;
	logic DTW_finish_r;
	
	logic similarity_word_r [0:499];
	logic [119:0] DTW_candidate_word_w [0:19], DTW_candidate_word_r [0:19];
	logic [119:0] DTW_word_r;
	logic [8:0] ptr_r, ptr_w;
	
	integer i;
	assign o_finish = finish_r;
	assign o_word = DTW_word_r;
	assign o_state = state_r;
	assign o_DTW_candidate_word = DTW_candidate_word_r;
	
	Similarity sim1(
		.i_similarity_clk(i_clk),
		.i_similarity_rst_n(i_rst_n),
		.i_similarity_start(similarity_start_r),
		.i_similarity_word(i_word),
		.o_similarity_finish(similarity_finish_r),
		.o_similarity_word(similarity_word_r)
	);
	
	DTW dtw1(
		.i_DTW_clk(i_clk),
		.i_DTW_rst_n(i_rst_n),
		.i_DTW_start(DTW_start_r),
		.i_DTW_word(i_word),
		.i_DTW_candidate_word(DTW_candidate_word_r),
		.o_DTW_finish(DTW_finish_r),
		.o_DTW_word(DTW_word_r),
		.o_state(DTW_state_r)
	);
	
	always_comb begin
		state_w = state_r;
		finish_w = finish_r;
		similarity_start_w = similarity_start_r;
		// similarity_finish_w = similarity_finish_r;
		DTW_start_w = DTW_start_r;
		// DTW_finish_w = DTW_finish_r;
		// DTW_word_w = DTW_word_r;
		// DTW_state_w = DTW_state_r;
		DTW_candidate_word_w = DTW_candidate_word_w;
		// similarity_word_w = similarity_word_r;
		ptr_w = ptr_r;
		
		case (state_r)
			S_IDLE: begin
				finish_w = 1'b0;
				if (i_start) begin
					similarity_start_w = i_start;
					state_w = S_CALC;
				end
			end
			S_CALC: begin
				similarity_start_w = 0;
				finish_w = DTW_finish_r;
				
				if (similarity_finish_r) begin;
					for (i = 0; i < DICT_SIZE; i = i + 1) begin
						if(similarity_word_r[i] == 1'b1) begin
							DTW_candidate_word_w[ptr_w] = dict[i];
							ptr_w = ptr_w + 1;
						end
					end
				end else if (pre_similarity_finish_r && !similarity_finish_r) begin
					DTW_start_w = 1'b1;
				end
				
				if (finish_r) begin
					state_w = S_DONE;
				end
			end
			S_DONE: begin
				finish_w = 1'b1;
				state_w = S_IDLE;
			end
		endcase
		
	end

	always_ff @ (posedge i_clk or posedge i_rst_n) begin
		if (i_rst_n) begin
			state_r                 <= S_IDLE;
			finish_r                <= 1'b0;
			similarity_start_r      <= 1'b0;
			// similarity_finish_r     <= 1'b0;
			pre_similarity_finish_r <= 1'b0;
			DTW_start_r             <= 1'b0;
			// DTW_finish_r            <= 1'b0;
			// DTW_word_r              <= 120'b0;
			DTW_candidate_word_r    <= '{20{120'b0}};
			// DTW_state_r             <= 3'b0; 
			// similarity_word_r       <= '{500{1'b0}};
			ptr_r                   <= 9'b0;

			
		end else begin
			state_r                 <= state_w;
			finish_r                <= finish_w;
			similarity_start_r      <= similarity_start_w;
			// similarity_finish_r     <= similarity_finish_w;
			pre_similarity_finish_r <= similarity_finish_r;
			DTW_start_r             <= DTW_start_w;
			// DTW_finish_r            <= DTW_finish_w;
			// DTW_word_r              <= DTW_word_w;
			DTW_candidate_word_r    <= DTW_candidate_word_w;
			// DTW_state_r             <= DTW_state_w;
			// similarity_word_r       <= similarity_word_w;
			ptr_r                   <= ptr_w;
		end
	end
endmodule

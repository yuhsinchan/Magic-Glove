module Dictionary (
    input          i_clk,
    input          i_rst_n,
    input          i_start,
    input  [119:0] i_word,
    output         o_finish,
    output [119:0] o_word,
    output [  1:0] o_state
    // output [119:0] o_DTW_candidate_word[0:19]
);
    parameter DICT_SIZE = 600;
    localparam bit [119:0] dict[0:DICT_SIZE - 1] = '{
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000110000000010100001110,
        120'b000000000000000000000000000000000000000000000000000000000001100100001100000101000000111000000101000000110000010100010010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010000110000010000000100100001010100010000,
        120'b000000000000000000000000000000000000000000000000000000000000111000000101000001010001010000010010000101010000111100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010000111100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010000110000000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000110000000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000001111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001000001010100010010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000010000010100000100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000000110001010100001100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000101000101100000010100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000010111000011110001001000000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100001110000000010000100000010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000101000100110000111100010000000100000001010100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000110000000100010000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000110010001010000010100000001010001001000010000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010000110000010000000011110000010100010000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011000000111100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100110000111100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000100000101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000111100010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000100000001010001000000010011000000010001001000000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000100110000110000000101,
        120'b000000000000000000000000000000000000000000000000000000000000000000010010000001010000100000010100000011110001001000000010,
        120'b000000000000000000000000000000000000000000001100000101010000011000010011000100110000010100000011000000110001010100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011110000111100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000100000011100000000100000010000100110001010100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000101000010110000000100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000001111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000101000001010000100000000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000010100001100,
        120'b000000000000000000000000000000000000000000000000000000000000000000010011000001010000100000010100000011110000110000000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000110001010100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100001011000000110001010100001100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000110000000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000101000011010000111100000011000011000000010100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011100000000100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010100010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000101000011010000111100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110001001000000101000010000001010000001111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000110000111000001111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100010010000011110001010000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100100000010100010110000001010000110000000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000100100000111100010000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110001001100001111000100100000001100000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000101000101100000010100001110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110000000100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100100000010100001000000101000000111100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000111100010010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000101000011100000111100000101000011010000111100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000011001000011000000110000000001000101000000111100010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000110010001010000001110000001010001011100010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010000110000000010000011010001010100001000,
        120'b000000000000000000000000000000000000000000000000000000000001001100010101000011110001001000001111000011010001010100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001100000100100000111100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001011000011110001000000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001010001001000000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011000000000100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010000001100001110000000010000100000000011,
        120'b000000000000000000000000000000000000000000000000000000000000010000001110000000010001001100010101000011110000100000010100,
        120'b000000000000000000000000000000000000000000000000000001000000010100001110000100100000010100000011000011100000111100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000011000000010001001000000111,
        120'b000000000000000000000000000000000000000000000000000000000001001100010011000001010000110000000101000100100000000100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010001100100000101,
        120'b000000000000000000000000000000000000000000000000000000000001001000000101000001110000000100001110000001010000010100010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001010000010100001011,
        120'b000000000000000000000000000000000000000000000000000000000000000000010010000001010000100000010100000011110000111000000001,
        120'b000000000000000000000000000000000000000000000000000100100000010100000111000100100001010100000010000011010000000100001000,
        120'b000000000000000000000000000000000000000000011001000100100001001000000101000000100001011100000001000100100001010000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100001011000011000000000100010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001100000010110000111000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000100110000000100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000100100000111100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100010111000011110000111000001011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000011000000010100000110,
        120'b000000000000000000000000000000000000000000000000000001000000010100010100000001010000110000010000000011010000111100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011100000001,
        120'b000000000000000000000000000000000000000000000000000000000001001000000101000001000000110000010101000011110000100000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000010100000100100000010100010011000100110000010100000100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100000011000000010000111000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000100000001010001100100001111000010100000111000000101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010100000101010001001000010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010001001100010101000000110001100000000101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000011010000000100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000100100000000100010000,
        120'b000000000000000000000000000000000000000000000000000000000000000000010011000011000000110000001111000100100001010000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001010100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100100000010100000110000001010001001000010000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010001011100001111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000011110001010000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100010011000001010001010100000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100010011000001010000110000000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000011100000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001100000101010000111100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100000011000001010000100000000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010001001000000011,
        120'b000000000000000000000000000000000000000000000000000000000001001100000101000001110000000100010011000100110000010100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000111100000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000001100000101010000010000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000100000011100000000100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011000000000100010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000101100000111100001100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000011000000000100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000001010000100000010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010000110000000100000011110000111100001110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000010000000111100001010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100000101000011100000111100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000011000011100001010100001100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000100000001010000010100001110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001010100000010,
        120'b000000000000000000000000000000000000000000000000000000000001010000010101000011100000100000000111000101010000111100000100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000101010000110000000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000000000100001111000100100000100000010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000101000011000000001000000001000100000000000100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000010011000001010000001100001110000000010000100000000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000100110000000100010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100100000010100000111000100100001010100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000001010000010100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010010000000010000010100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000010100000100110000010100010100000011100000111100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000010110000000100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000010000010100001010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010000011100001110000000010001001000001111,
        120'b000000000000000000000000000000000000000000000000000000000000000000010100000011100000010100000100000101010001010000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000001010000010100000110,
        120'b000000000000000000000000000000000000000000000000000000000000110000001100000000010000001000010100000011110000111100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000100000100100000111100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000010110000111100001010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000100110000111100001100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000100100000010100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000111100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000010000010100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000011000000000100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011000000000100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000101010000100000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000010010000001010000010000001110000001010000110000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000001100001110000101010001001000000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010100000100110000000100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000111000101010000111100000011,
        120'b000000000000000000000000000000000000000000000000000000000001100100000001000001000001001000010101000101000000000100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010000111000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000111000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010101000011110000001000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010001001100000001000001010000110000010000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001100000011110000100000010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000011000000010100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100100000010100010000000100000001010100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000001010000010100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000010000010100011001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100010000000001010001010000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000111100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000000010100000111000100100000111100000110,
        120'b000000000000000000000000000000000000000000000000000011000001010100000110000100100000010100000100000011100000111100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001010100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000100100000111100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000111100001110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100100000010100000011000011100000000100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000110010000110000000101000011100000111100001100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001110000101010000111100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011110000111100000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011000110010000000100000100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000011000000111000001111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000101110000111100010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001110000011110000110100000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000011001000100000001000000000001000010000000111000010101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011000001010000011100000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000001100000011110001001000010100000011100000111100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000010000010100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000001001000001111000001100000011000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010100001100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011000000111100000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000101000101010001001000000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000001010000001100000000010000010100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000101010000111100011001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000110010000101100000001000001010000111000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000110010000110000000100000000010000010100000100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010000000000010001001000000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000101000001110000111000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000000100000000111000101010000000100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000110010000001000000010000101010000100000000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000100100000111100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000010000010100001110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010001001000001111000001100000010100000010,
        120'b000000000000000000000000000000000001001000000101000010000001010000000001000001100000010000001110000000010001001000000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000100110000000100000101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100110000010100010010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000011110000111100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110000111100001110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000010101000011110001001000010000,
        120'b000000000000000000000000000000000000000000000000000000000000000000010010000001010001011000001111000000110000010100010010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000101000001000000110000000101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010001001000010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100110000010100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000001100000101010000011000000101000100100000000100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000100000010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000010011000011100001001000010101000101000000010100010010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110001010100010000000011010000000100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000010011000011010000111100010100000101000000111100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000100100000010100010110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100110001010100001010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110000111100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100001100000100000000010100010010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000100000001010000011100010010000000010000100000000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001010001001100010101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000101000101000000111000000101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000011100000101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111000011110000100000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000101000001010001001000000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011000000111100000100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000111100010100,
        120'b000000000000000000000000000000000000000000000000000000000000010000000101000101000000000100000101000001100000010100000100,
        120'b000000000000000000000000000000000000000000000000000000000001001000000101000001110000111000000001000100100001010000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000101010000111100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000110000000100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100000001000001010001000000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000001000000000101000000110001100000000101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010011000100100000111100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000011000101010000111100010100,
        120'b000000000000000000000000000000000000000000000000000000000000111000001111000100110000010000001110000000010001001000000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100100000010100001100000011000000000100010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000011100000010100010110000001010000110000000101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000001001100000101000101000000000100001100,
        120'b000000000000000000000000000000000000000000000000000000000000000000010010000001010000100000010100000000010000010100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000101000000111100000010,
        120'b000000000000000000000000000000000000000000000000000001010001010000000001000011000000111100000011000011110000100000000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000101000101110000111100010000,
        120'b000000000000000000000000000000000000000000000000000000000001001000000101000011010000111100010100000100110001010100000011,
        120'b000000000000000000000000000000000001001100001110000011110000110000000101000011010001001000000101000101000000000100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011000001010001011100001111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000100100001010100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000000010001010000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100001011000000110000000100001100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000100000001010000110000001100000001010000110100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000010101000001100001011100000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010010000000010000110100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011000001010100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010110000000010000010100001100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000001000000000100001100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000101110000111100000100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100100000111100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000100100001010100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000010000010100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110001010100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000101010001001000010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000001110000101010000111100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000011100000010100000100000100100000000100000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010010000001010000100000010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010000000100000100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000001001100000101000001000000111100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010100000101010000111100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000000010100010010000001110000010100010010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011000100110000000100010000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000000010001001000000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100100000010100001100000011110000111100000011,
        120'b000000000000000000000000000000000000000000000000000011100000000100001101000001010000110000010100000011100000010100000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010000000100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000110000011000000010100010011000100100000010100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100000011000000010000110000000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010101,
        120'b000000000000000000000000000000000000000000000000000001000000010100010100000100110000010100000111000001110001010100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000101100000111100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110000000100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000000100000011,
        120'b000000000000000000000000000000000000000000001110000011110000110000000101000011010001001000000101000101000000000100010111,
        120'b000000000000000000000000000000000000000000010100000011100000000100010010000101010000000100010100000100110000010100010010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001010100000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010010000011110000100000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000001000001010001001000000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100100001010100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100100000010100010100000100110000000100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010001001000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000010100000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000001010000010100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000101000101000000011000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110000010000001110000101010000111100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110001100100000001000101110000110000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000101000100110001010100000001000000110000010100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000100000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000010000101010000111100000100,
        120'b000000000000000000000000000000000000010100001000000000110000000100001000000000110000000100001101000011110001010000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011000100100000000100000101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100100000010100010111000100110000111000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000001001100000101000011100000111100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000111000001111000000110000010100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001010100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100000100000011100000000100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000011100000000100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000001000000111100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001010100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000010000000011110000110000000101000101100000010100000100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000011000000000100010000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010110001001100000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000011100000111100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000110010000110000000101000101100000111100001100,
        120'b000000000000000000000000000000000000000000000000000101000001001100000001000001100000101100000001000001010001001000000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110000101100000011000011110000111000001011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000110010001010000001110000001010000110000010000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000010100010000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010011000011100000010100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000011001000010000001010000001100000000010000010100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000001010001011000001111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000010000111000000001000011100000000100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000111000011100000000100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010001001000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000101000100100000100000010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000011010000000100000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000100100000000100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000011001000101000000111000000101000101100000010100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000101000011100001011100001111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100010000000100000000000100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000110010000110000000100000100100000000100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000101000011110000100000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100110000111100001100,
        120'b000000000000000000000000000000000000000000000000000000000000010100001000000000110000000100000100000000010000010100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000101000010110001001100000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000010000100000010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010000100000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000100000001010000111000010111000011110001001000000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000101010000111100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000010100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000001110000001010000010100010111000101000000010100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000011100000010100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000101010000111100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100100000010100001000000101000000000100010010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000111100000100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000011110000100000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000101110000111100001100000011000000010100011001,
        120'b000000000000000000000000000000000000000000000000000000000000000000011001000101000000100000000111000101010000000100001110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010100000101010000111100011001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000011110001001000000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000001110000111000001111000100100001010000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010000100000010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000111100011001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000110000001111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011000000000100000011,
        120'b000000000000000000000000000000000000000000000101000011000000001000000001000010110001001000000001000011010000010100010010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000111100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110000010100001011000011110000110100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001011100001111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100100000010100011001000101110000000100001100,
        120'b000000000000000000000000000000000000000000000000000110010000000100000100000100100000010100010100000100110000010100011001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000010100010011000101010000000100010000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011000000111100010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011000001010001100100000101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000100110000000100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100001100000001000000000100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010010000000010000010100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011000000010100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000000111000000101000100100000000100010000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000001000001010001001000010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000100000010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111000011110000110000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011110000111100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000001010001001000000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000100100000111100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000101000010110000000100010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000101000001010000110000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000010100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000010011000101010000111100010110000100100000010100001110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000000100000000100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001000000000100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010011000011110000100000010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000011000000000100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100100000010100010100000100110000000100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110000000100001100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000100100000111100011001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000111100000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010100010010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001110000011110000110000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100001100000011000000000100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000011010000111100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000111000100100000000100001100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000000101000001000000111000010101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000010100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100100000010100010100000101000000010100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000110000010101000011110000100000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000010100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000110010000110000001100000000010000010100010010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000011110000111100010000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000011110001010000000001000011010000111100010100,
        120'b000000000000000000000000000000000000000000000101000011000000001000000001000011100000111100010011000000010000010100010010,
        120'b000000000000000000000000000000000000000000000000000001010000011100000100000001010000110000010111000011110000111000001011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000101000100100000111100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000101000000000100010000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000100010010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000011000000010100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010001001100010010000101010000111100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110000101100001110000000010000100000010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010001001100010101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010110000000010001001000000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000101000001010001010100010001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000100110001010100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110000010100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000010100011001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100001110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000110010000000100000100000011100001010100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010011000101010000111100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100001110000011100001010100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010000110000010000000101010000111100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001010000010100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000010011000100100000000100000101000100000001000000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100100000010100001110000100100000111100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000001010000100000010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010011000001010000100000010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011000001010000111100000100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111000011110001001000000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000010011000001000000111000000101000100000000010100000100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000010110000000100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001010000010100001110,
        120'b000000000000000000000000000000000000000000000000000001000000010100010100000100110001010100000001000010000001100000000101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100001011000011110000111100001100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000100110000111100001110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100110000111100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000111000010101000011110001001000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000110000001100000111100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000101100000000100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100110000000100001100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001011100001111000011000000110000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011000100110000111100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100000001000001010001010000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100001100000001010000010100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001110000011110001001000010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011000000010100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000001100000101010000000100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100001010100001111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000100000001010001001000000100000011100001010100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000011000000111100001111000010000000001100010011,
        120'b000000000000000000010010000001010001010000001000000001110001010100000001000001000000010000001110000000010001001000000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000101000001010100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000000110000000100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000011100000111100010011000100100000010100010000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000000110000010100001110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100010100000100100000111100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000011110000111100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100001011000011000000000100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000100000011110000111100000110000000010000010100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100000011000011100000000100001110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000100100000010100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100010100000100100000000100010000,
        120'b000000000000000000000000000000000001001000000101000010000001010000001111000011010000010000001110000000010001001000000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100010010000001110000111000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010011000011000000000100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000111100001110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000001010000100000010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000110000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000101000000000100001100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001010100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000001111000011010000010100001100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000101000001110000111000000001000100100001001000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000101000100100000011100000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100010010000100100001010100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010100000000010000010100000100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010010000001010000100000010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000101000011000000001000010101000011110001001000010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000010000010100001110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001100000101010000111100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010010000000010001010000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010011000001010001010100000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011110000111100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010011000101010001001000010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001100000001010000110100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100001111000010100000111000000101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000001111000101100000000100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000011010001010100000100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000100000100100000000100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100000001000001010001001000000100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000011000000111100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011100000000100010111,
        120'b000000000000000000000000000000000000000000000000000000000000010000000101000011100000010100010000000100000000000100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111000011110000111000001011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000010100001011000011000000000100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000010011000001010000111000001111000001110001100100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001100000000010000100000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000010100010110000100100000010100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110000010100001110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110000110000000001000101010001000100000101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000010000010100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001100000100000001000000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000010000010100000100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000010000100000010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000010110000000100010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011000000111100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000011010000111100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000010100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001110000101010000111100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000000100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000011100000010100010100000100110000000100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001110000000010000110000010000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010000010100010010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100000100000000010000010100010010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100001101000001010000010100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000010000100000010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001010100001111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100010010000100100000111100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000111000001111000110010000010100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001000001010000100000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010000000100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001010000111000001011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001100000000110000111000010101,
        120'b000000000000000000000000000000000000000000000000000000000000000000001101000001010000110000000010000011110001001000010000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010110000011110000001000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000010000010100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000000010001011100000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010000000100001101,
        120'b000000000000000000000000000000000000000000000000000000000000011000001100000001010001001100010010000101010000111100011001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000001000000000101000000110000001100000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000011000101000000000100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000100000001010000010000001110000101010000111100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000001000011010000111100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000001000100000000000100001010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010010000000010000100000010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011000001111,
        120'b000000000000000000000000000000000000000000000000000000000001100100000001000001000001100100010010000001010001011000000101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000011000011100000000100000100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000011100000111100001110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000000010000110000010000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001101000101010000100000010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000010100001100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000110010001001000001111000011010000010100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000111000001111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000100,
        120'b000000000000000000000000000000000000000000000000000000000001001000000101000101000000100000000111000101010000000100000100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011000000010100010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000011100000111100001100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000110010000010000000101000001010001001000000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001011000011110001001000000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000000010100000101000100100001010000010011,
        120'b000000000000000000000000000000000000000000000000000000000001011100001111000100100001001000001111000011010000111100010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000100000001010001001100010011000001010001001000000100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000001010000100000010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100010010000100100000111100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000101110000111100001100000011000000010100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000101010000111100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000010000111100000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010001001100000101000001010000100000000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110000000100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100010010000100100000000100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000010110000000100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000011100000010100001011000011110001001000000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000001111000011010001010100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000011110000111100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001011100001111000011000000010100000010,
        120'b000000000000000000000000000000000000000000000000000000000000000000010011000100100000010100010111000100110000111000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000011100000111100010011000000010000010100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000001111000011010001010100010010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000010100010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001110000011110000110000000001,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110001010100001111000011010000000100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010001010100000111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000111100001010,
        120'b000000000000000000000000000000000000000000000000000000000000000000010010000001010000111000010100000100100000000100010000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000100100000010100001000000101000000000100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000011110000111100001100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100110000000100000101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011000000010100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000101000101100000010100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011000000010000010100010111,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011000000000100001000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100000001000001000000111100010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000001100000110000000101000100110001100100001101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111000001010000111000001011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100010010000001010001011000000101,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000001111000011000000111100000011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000000010000010100010000,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100010010000101010000111100011001,
        120'b000000000000000000000000000000000000000000000000000000000000000000010011000101010000111100001100000000010000010100001010,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000011010000111100010011,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000101110000111100001100000011000000111100000110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000010101000011110000110000000110,
        120'b000000000000000000000000000000000000000000001100000101010000011000010100000010000000011100010101000011110000100000010100,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000011010000000100001110,
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100001001
    };

    localparam S_IDLE = 3'd0;
    localparam S_IREV = 3'd1;
    localparam S_CALC = 3'd2;
    localparam S_OREV = 3'd3;
    localparam S_DONE = 3'd4;

    logic [2:0] state_r, state_w;
    logic finish_r, finish_w;

    logic [119:0] i_reverse_word_w, i_reverse_word_r, o_reverse_word_w, o_reverse_word_r, tmp_word_r, tmp_word_w;
    logic [4:0] i_word_length, o_word_length;
    logic [4:0] counter_r, counter_w;

    logic similarity_start_r, similarity_start_w;
    logic similarity_finish_r, pre_similarity_finish_r;
    logic similarity_finish;
    logic [2:0] DTW_state_r;  // debug
    logic DTW_start_r, DTW_start_w;
    logic DTW_finish_r;

    logic [9:0] similarity_word_r[0:19];
    logic [119:0] DTW_candidate_word_w[0:19], DTW_candidate_word_r[0:19];
    logic [119:0] DTW_word_r;
    logic [8:0] ptr_r, ptr_w;

    integer i;
    assign o_finish = finish_r;
    assign o_word = o_reverse_word_r;
    assign o_state = state_r;
    // assign o_DTW_candidate_word = DTW_candidate_word_r;
    assign i_word_length = (i_word[7:0] != 8'b0) + (i_word[15:8] != 8'b0) + (i_word[23:16] != 8'b0) + (i_word[31:24] != 8'b0) + (i_word[39:32] != 8'b0) + (i_word[47:40] != 8'b0) + (i_word[55:48] != 8'b0) + (i_word[63:56] != 8'b0) + (i_word[71:64] != 8'b0) + (i_word[79:72] != 8'b0) + (i_word[87:80] != 8'b0) + (i_word[95:88] != 8'b0) + (i_word[103:96] != 8'b0) + (i_word[111:104] != 8'b0) + (i_word[119:112] != 8'b0);
    assign o_word_length = (DTW_word_r[7:0] != 8'b0) + (DTW_word_r[15:8] != 8'b0) + (DTW_word_r[23:16] != 8'b0) + (DTW_word_r[31:24] != 8'b0) + (DTW_word_r[39:32] != 8'b0) + (DTW_word_r[47:40] != 8'b0) + (DTW_word_r[55:48] != 8'b0) + (DTW_word_r[63:56] != 8'b0) + (DTW_word_r[71:64] != 8'b0) + (DTW_word_r[79:72] != 8'b0) + (DTW_word_r[87:80] != 8'b0) + (DTW_word_r[95:88] != 8'b0) + (DTW_word_r[103:96] != 8'b0) + (DTW_word_r[111:104] != 8'b0) + (DTW_word_r[119:112] != 8'b0);

    Similarity sim1 (
        .i_similarity_clk(i_clk),
        .i_similarity_rst_n(i_rst_n),
        .i_similarity_start(similarity_start_r),
        .i_similarity_word(i_reverse_word_r),
        .o_similarity_finish(similarity_finish_r),
        .o_similarity_word(similarity_word_r)
    );

    DTW dtw1 (
        .i_DTW_clk(i_clk),
        .i_DTW_rst_n(i_rst_n),
        .i_DTW_start(DTW_start_r),
        .i_DTW_word(i_reverse_word_r),
        .i_DTW_candidate_word(DTW_candidate_word_r),
        .o_DTW_finish(DTW_finish_r),
        .o_DTW_word(DTW_word_r),
        .o_state(DTW_state_r)
    );

    always_comb begin
        state_w = state_r;
        finish_w = finish_r;
        similarity_start_w = similarity_start_r;
        // similarity_finish_w = similarity_finish_r;
        DTW_start_w = DTW_start_r;
        // DTW_finish_w = DTW_finish_r;
        // DTW_word_w = DTW_word_r;
        // DTW_state_w = DTW_state_r;
        DTW_candidate_word_w = DTW_candidate_word_w;
        // similarity_word_w = similarity_word_r;
        ptr_w = ptr_r;

        i_reverse_word_w = i_reverse_word_r;
        o_reverse_word_w = o_reverse_word_r;
        counter_w = counter_r;
        tmp_word_w = tmp_word_r;

        case (state_r)
            S_IDLE: begin
                finish_w = 1'b0;
                if (i_start) begin
                    state_w = S_IREV;
                    counter_w = 0;
                    tmp_word_w = i_word;
                end
            end
            S_IREV: begin
                if (counter_r < i_word_length) begin
                    i_reverse_word_w = {i_reverse_word_r[111:0], tmp_word_r[7:0]};
                    tmp_word_w = tmp_word_r >> 8;
                    counter_w = counter_r + 1;
                end else begin
                    state_w = S_CALC;
                    similarity_start_w = 1'b1;
                    counter_w = 0;
                end
            end
            S_CALC: begin
                similarity_start_w = 0;

                if (similarity_finish_r) begin
                    for (i = 0; i < 20; i = i + 1) begin
                        DTW_candidate_word_w[i] = dict[similarity_word_r[i]];
                    end
                end else if (pre_similarity_finish_r && !similarity_finish_r) begin
                    DTW_start_w = 1'b1;
                end

                if (DTW_finish_r) begin
                    state_w = S_OREV;
                    counter_w = 0;
                    tmp_word_w = DTW_word_r;
                end
            end
            S_OREV: begin
                if (counter_r < o_word_length) begin
                    o_reverse_word_w = {o_reverse_word_r[111:0], tmp_word_r[7:0]};
                    tmp_word_w = tmp_word_r >> 8;
                    counter_w = counter_r + 1;
                end else begin
                    state_w = S_DONE;
                    counter_w = 0;
                end
            end
            S_DONE: begin
                finish_w = 1'b1;
                state_w  = S_IDLE;
            end
        endcase

    end

    always_ff @(posedge i_clk or posedge i_rst_n) begin
        if (i_rst_n) begin
            state_r                 <= S_IDLE;
            finish_r                <= 1'b0;
            similarity_start_r      <= 1'b0;
            // similarity_finish_r     <= 1'b0;
            pre_similarity_finish_r <= 1'b0;
            DTW_start_r             <= 1'b0;
            // DTW_finish_r            <= 1'b0;
            // DTW_word_r              <= 120'b0;
            DTW_candidate_word_r    <= '{20{120'b0}};
            // DTW_state_r             <= 3'b0; 
            // similarity_word_r       <= '{500{1'b0}};
            ptr_r                   <= 9'b0;
            i_reverse_word_r <= 120'b0;
            o_reverse_word_r <= 120'b0;
            tmp_word_r <= 120'b0;
            counter_r <= 4'b0;

        end else begin
            state_r                 <= state_w;
            finish_r                <= finish_w;
            similarity_start_r      <= similarity_start_w;
            // similarity_finish_r     <= similarity_finish_w;
            pre_similarity_finish_r <= similarity_finish_r;
            DTW_start_r             <= DTW_start_w;
            // DTW_finish_r            <= DTW_finish_w;
            // DTW_word_r              <= DTW_word_w;
            DTW_candidate_word_r    <= DTW_candidate_word_w;
            // DTW_state_r             <= DTW_state_w;
            // similarity_word_r       <= similarity_word_w;
            ptr_r                   <= ptr_w;
            i_reverse_word_r <= i_reverse_word_w;
            o_reverse_word_r <= o_reverse_word_w;
            tmp_word_r <= tmp_word_w;
            counter_r <= counter_w;
        end
    end
endmodule

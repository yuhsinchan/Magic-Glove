module Pseudo_random (
    input i_reset,
    input [3:0] i_seed,
    input i_jingyuanhaochiang,
    output [3:0] o_lfsr_random, 
);

endmodule
module similarity(
	input i_similarity_clk,
	input i_similarity_rst_n,
	input i_similarity_start,
	input [119:0] i_similarity_word,
	output o_similarity_finish,
	output o_similarity_word[0:499],
);

	parameter COUNT_DICT_SIZE = 500;
	localparam bit [103:0] count_dict[0:COUNT_DICT_SIZE - 1] = '{
		120'b00000000000000010000000000000000000100000000000100000000000000000000000000000000000000000001000000000000,
		120'b00000000000000000000000000010000000000000000000000000000000000000000000000010000000000010000000000000000,
		120'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000100000000000000000000,
		120'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000001,
		120'b00000000000000000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001,
		120'b00000000000000000000000000000000000000000000000000010000000000000000000100000000000000000000000000000000,
		120'b00000000000000000000000000000000000100000000000100000000000000000000000000000000000100000000000000000000,
		120'b00000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000000001,
		120'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000,
		120'b00000000000000000000000000010001000000000000000000000000000000000000000100010000000000000000000000000000,
		120'b00000000000000010000000000010000000000000000000000000000000000000000000100010000000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000,
		120'b00000001000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000,
		120'b00000000000000000000000000010000000000000000000100010000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000,
		120'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000001,
		120'b00000000000000000000000000000000000100000000000100000001000000000000000000000000000100000000000000000000,
		120'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000001,
		120'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001,
		120'b00000001000000000000000100000000000100000000000100000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001,
		120'b00000000000000000001000000000000000000000000000000000000000000000000000000010000000000010000000000000001,
		120'b00000000000000010000000000000000000000000000000000010000000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000000000000000100000000000100000001000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001,
		120'b00000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000001,
		120'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000,
		120'b00000000000000010000000000000000000000000000000000000000001000000000000100000000000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000100000001000000000000000000010000000000010000000000000000,
		120'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000001,
		120'b00000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000100010000000000000000000100000000000000000000000000000000000000000000000000010001,
		120'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000,
		120'b00000000000000000000000000000000000000000001000000000000000000000000000000000001000000010000000000000001,
		120'b00000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000001,
		120'b00000000000000000000000000000001000100000000000000000000000000000000000000010000000000010000000100000001,
		120'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000100100000000000000000,
		120'b00000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000010000,
		120'b00000000000000000000000100000000000100000000000100000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000100010000000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000000010000000100000000000100000000000000000000000000010000000000010000000000000000,
		120'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001000000000000,
		120'b00000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000010000000100000000001000100001000000000000001000000000000100000000000000000001,
		120'b00000000000000000000000000010000000000000000000000000001000000000000000100000000000000010000000000000000,
		120'b00000001000000000000000000010000000000000000000000000000000000000000000000010000000000010000000000000000,
		120'b00000000000000000000000000010001000000000000000000000000000000000000000100000000000000010000000000000000,
		120'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000,
		120'b00000000000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000,
		120'b00000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001,
		120'b00000000000000010000000000010000000000000000000000000000000000000000000000010000000000000000000000000001,
		120'b00000000000000010000000000000000000000000000000000000000000000000000000100100000000000000000000100000000,
		120'b00000000000000000000000000010000000100000000000000000000000000000000000100010000000000010000000000000000,
		120'b00000000000000010000000000000001000000000000000000010000000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000100010000000000000000000100000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000100000001000000000000000000000000000000000000000000000000000000010000000000000000,
		120'b00000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001,
		120'b00000000000000000000000000010000000100000000000000000000000000000000000000010000000000100000000000000000,
		120'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000100000000000000000,
		120'b00000001000000000000000000000000000000000000000100010000000100000000000000000000000000000000000000000000,
		120'b00000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000000001000000000000000000000000000000000000000100010000000000000000000000000000,
		120'b00000000000000010000000000000000000000000000000000010000000000000000000000010000000000010000000000000000,
		120'b00000000000000000000000000100000000000000000000100010000000000000000000000000000000000000000001000000001,
		120'b00000000000000000000000000000000000100000000000000000000000000000000000000010000000000100000000000000000,
		120'b00000000000000000000000100000011000000000000000000010000000000000000000100000000000000010000000000010000,
		120'b00000000000000010000000000000000000000000000000100000000000000000000000000010000000000000000000000000000,
		120'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000010000,
		120'b00000000000000000000000000000001000000000000000100000000000100000000000000000000000000000000000000000001,
		120'b00000000000000010000000000000000000000000000000100010000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000000000000000000001000000000000000100000000000000010000000000010000000000000000,
		120'b00000000000000000000000000010000000000000000000000000000000000000000000000000001000000010000000000000000,
		120'b00000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000000000,
		120'b00000000000000010001000000000000000000000000000000000000000000000000000100000000000000010000000000000000,
		120'b00000000000000000000000000000000000000000000000100100000000100000000000100000000000000010000000000000000,
		120'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000,
		120'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000000010001000100000000000000000000000000000000000100000000000100000000000000000000,
		120'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001,
		120'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000100000000000010000,
		120'b00000000000000010000000100000000000000000000000100000000000100000000000000000000000000000001000000000000,
		120'b00000000000000010000000000000000000000000000000100000000000000000000000000010000000000000000000000000000,
		120'b00000000000000010000000000000000000100000000000000000000000000000000000000000000000000100000000000000000,
		120'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000001000000000010000100000000000000000000000000000000000100000000000000100000000100000000,
		120'b00000000000000000000000000000001000000000000000100000001000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000000010001000000000000000000000000000000000000000000010000000000100000000000000000,
		120'b00000000000000000000000000000000000000000000000000000000000100010000000100000000000000000000001000000000,
		120'b00000000000000000000000000010001000000000000000000000000000000000000000100000000000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000000000000000100010000000100000000000000010000000000000000,
		120'b00000000000000000001000000000001000100000000000000000000000000000000000100000000000000100000000100000000,
		120'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000010000000000000000000000010000000000000000000000010000000000000000000000000001,
		120'b00000000000000000000000000000000000000000000000000010000000000000000000100000000000100000001000000000000,
		120'b00000000000000000000000000000000000100000001000000000000000000000000000100000000000000010000000100000000,
		120'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000010001000000000001,
		120'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001,
		120'b00000000000000000000000000010000000000000001000100000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000000000000000000010000100000000000100000000000000000000000000100000000000000000,
		120'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000001,
		120'b00000000000000000000000000010001000000000000000000000000000100000000000100000000000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000000010001000000000000000000000000000000010000000000000001,
		120'b00000000000000000000000100010001000000000000000000000000000000000001000000000000000000000000000000000000,
		120'b00000000000000000001000000000000000100000000000100000000000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000000100001000000000000000000000000000000000000000000000000000000010000000000000001,
		120'b00000001000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000001,
		120'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001,
		120'b00000000000000000000000000010000000000000000000100010000000000000000000100000000000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000000000001000100000000000100000000000000010000000000000001,
		120'b00000000000000010000000000010000000000000000000100000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000010000000000000000000000000000000100000000000000100000000000010000000000000001,
		120'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000,
		120'b00000000000000010000000000000000000100000000000100000000000100000000000000000000000000000001000000000000,
		120'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000,
		120'b00000000000100000000000000010000000000000000000000010000000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000100000001000000000000000000000000000000000000000000000000000000010001000000000000,
		120'b00000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000,
		120'b00000000000000010000000000000000000100000000000100000000000000010000000000000000000000000000000000000000,
		120'b00000000000000000000000000010001000000000000000000000000000100000000000000000000000000000000000000000001,
		120'b00000000000000000000000000010001000000000000000100000001000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000100010001000100000001000100000000000000000000000000000000000000000001000100000000,
		120'b00000000000000000000000100000001000000000000000000000001000000000000000100000000000000000000000100000000,
		120'b00000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000,
		120'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000010,
		120'b00000000000000000000000000000000000000000000000000000001000000010000000000000000000000010000000000000001,
		120'b00000000000000000000000000010000000000000000000000000001000000000000000000010000000000010000000000000000,
		120'b00000000000000000000000100000001000000000000000100000000000100000000000000010000000000000001000000000000,
		120'b00000000000000000000000100010000000100000001000100000000000000000000000000000000000000000001000100000000,
		120'b00000001000000000000000000010010000000000000000000000001000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000000010001000000000001000100000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000000000000100000000000000000000000000000000000000010000000000010000000000000000,
		120'b00000001000000000000000000010000000000000000000000000000000000000000000100000000000000000000000100000000,
		120'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000001,
		120'b00000001000000000000000000000000000000000001000100000000000100000000000100000000000000000000000100000000,
		120'b00000000000000000000000100000000000100000000000000010001000000000000000000000000000000010000000000010000,
		120'b00000000000000000000000100000001000000000000000000000000000000000000000000010000000000000000000100000000,
		120'b00000000000000000000000000000001000000000001000000000000000100000000000000000000000000100000000000000001,
		120'b00000000000000000001000000000000000000000000000000000000001000000000000100000000000000010000000000010011,
		120'b00000001000000000000000000010000000100000001000100000000000000000000000100010001000000000000000100000000,
		120'b00000000000000000000000100010001000100000010000100000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000000010000000000000000000000001000000000000000000000001000000100000000000000001,
		120'b00000000000000000000000000010000000100000000000000000000000000000000000000000000000100010000000000000001,
		120'b00000000000000000000000000010001000000000000000000000000000000000000000000000000000000010000000000010000,
		120'b00000000000000010000000000010001000100000000000100000000000000000000000000000000000100010000000000000001,
		120'b00000000000000000000000000010000000000000000000000010000000000000000000000010000000000010000000000000000,
		120'b00000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000001,
		120'b00000000000000000000000000000000000000000000001000000000000000000000000000000001000000000001000000000000,
		120'b00000000000000000001000000000000000000000000000100000000000000000000000100000000000000010001000000000000,
		120'b00000000000000010000000000000000000000000000000000000000001000000000000000000000000000010000000000000000,
		120'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000,
		120'b00000000000000010000000000000000000100000000000000000000000000000000000000010000000000100000000000000000,
		120'b00000000000000000000000000000000000000000000000100010000000000000000000100000000000100000000000000000000,
		120'b00000000000000000000000000010001000100000000000000000000000000000000000100010001000000000000000000000000,
		120'b00000000000000000000000100000000000000000001000000000000000100000000000100000000000000000000000100010000,
		120'b00000000000000000000000000000001000000000000001000000000000000010000000000000000000000000000000000010000,
		120'b00000000000000000000000000000000000000000000000000000000000000000000000100100001000000000000000000000000,
		120'b00000000000000000000000000000001000000000000001000000000000100000000000000010000000000000000000100000000,
		120'b00000000000000000000000100010000000100000000000100000000000000000000000000100001000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000100000001,
		120'b00000000000000000000000000000001000000000000000000010000000100010000000100000000000000000000000000000000,
		120'b00000000000000000000000000000001000000000000000000000000000000000000000000010000000000010000000000000000,
		120'b00000000000000010001000000000000000100000000000000000000000000000000000100000000000000100000000000000000,
		120'b00000001000000000000000000000001000100000000000000000000000000000000000000000000000000010000000000000001,
		120'b00000000000000000000000000000000001000000000000100000000000000000000000000000000000000010001000000000000,
		120'b00000001000000000001000000000000000100000000000000000000000000000000000000000000000000010000000000000000,
		120'b00000001000000000001000000000000000100000001000000000000000000000000000100000000000000000000000100000001,
		120'b00000000000000000000000000000000000000000000001000000000000000010000000000000000000000000000000000010000,
		120'b00000000000000000000000000010001000000000000000000000001000000000000000100000000000000010000000000000000,
		120'b00000001000000000000000000000000000000000001000100010001000000000000000000000000000000000000000100000001,
		120'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000010001000000000001,
		120'b00000000000000000000000100000000000100000001000100000000000000000000000000000001000000000000000000000000,
		120'b00000000000100000000000000000001000000000000000000000000000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000100001000000000000,
		120'b00000001000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000001,
		120'b00000000000000000000000100000001000100000000000000000000000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000000000001000000000000000000000000000000000000000100000000000000000001000000000001,
		120'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000,
		120'b00000000000000000000000000000001000000000000000100000000000000000000000000000000000000010001000000000000,
		120'b00000000000000000000000000010001000000000000000000000000000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000100000000000100000000000000010000000000000000000000000000000000010001000000000000,
		120'b00000000000000000000000000000000000100000000000000010000000100000000000000000001000000100000000000000001,
		120'b00000000000000000000000000000001001000000000000000000000000000000000000000010000000000100000000100000001,
		120'b00000001000000000001000100010001000100000000000000010000000000000000001000000000000000010000000000000000,
		120'b00000001000000000000000100000000000100000000000000010000000000000001000000000000000000000000000000000010,
		120'b00000000000000000000000000000000000000000000000000000001000100000000000100000000000000000000000000000001,
		120'b00000000000000000000000100000000000000000000000000000000001000000000000000000000000100000000000000000000,
		120'b00000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000000001,
		120'b00000000000000010001000000000001000100000000000000000000000000000000000100000000000000100000000000000000,
		120'b00000000000000000000000000000000001000000001000100000001000000000000000000000001000000000000000000000001,
		120'b00000000000000000000000000000000000000000000000000000000000100000000000100000000000100010000000000000000,
		120'b00000000000000010000000000000000000000000000000100010000000000010000000000000000000000000000000000000000,
		120'b00000000000000000000000000000001000000000000000000000001000000000000000000000001000000010000000000000001,
		120'b00000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001,
		120'b00000001000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000001,
		120'b00000000000000000000000000010000000000000000000000100010000000000000000000000001000000100000000000000010,
		120'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000010000000100000001000000000000000000000000000000000000000000000000000000000001,
		120'b00000000000000000000000100000000000000000000000100000000000100000000000000000000000000000001000100000000,
		120'b00000000000000000000000000010000000100000000000000000000000000000000000000000001000000010000000000000001,
		120'b00000000000000000000000100010000000000000000000000010000000000000000000100000000000000010001000000000000,
		120'b00000000000000000000000000010000000000000000000100000000000100000000000000010000000000010000000000000000,
		120'b00000000000000000000000000000000000100000000000000000000000100000000000000000000000000010000000000000001,
		120'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000,
		120'b00000000000000000000000000010000000000000000000000000001000000000000000100000000000000010000000000000000,
		120'b00000000000000000000000000100000000100000000000100110000000100000000001000000000000000010000000000000010,
		120'b00000000000000000000000000010000000100000000000000010000000000000000000000000000000000100000000100000000,
		120'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010001,
		120'b00000000000000000000000100010001000000000000000000000001000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000010001000100000000000100000000000000000000000000000000000000010000000000000000,
		120'b00000000000000000001000000010000000100000000000000000000000100000000000000000000000000010000000000000001,
		120'b00000000000000000000000000010001000000000000000100010010000000000000000000000000000000010000000100000000,
		120'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000010001000000000001,
		120'b00000000000000000001000000010000000000000001000100010001000100000000000000000000000000110001000000000000,
		120'b00000000000000000000000000010000001000000001000100000000000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000000000000000000000000000100000000000000000000000000000000001000000000000000000000,
		120'b00000000000000000000000000000000000100000000000000000010000000000000000000000000000000100000000000010000,
		120'b00000000000000000000000000010001000000000000000000000000000100000000000100000000000000010001000000000001,
		120'b00000000000000000000000000000000000000000000000000010000000100000000000100000000000000010000000000000000,
		120'b00000000000000000000000000010001000100000000000000000001000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000000000000000100000000000100000000000000000000000000000000000100100000000000010000,
		120'b00000000000000000000000000010001000000000000000100000000000100000000000000010000000000010000000000000000,
		120'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000000000,
		120'b00000000000000000000000000000001000000000000000000010000000000000000000000000000000000010001000000000000,
		120'b00000000000000000000000000010000000100000000000000000000000000000000000100010001000000000000000000000000,
		120'b00000001000000000000000000010000000000000001000000000000000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000100000001000000000000000000000000000000000000000000000000000000100000000100010001,
		120'b00000000000000000000000000000000000000000000000100000000001000000000000000000000000000000000000100000001,
		120'b00000000000000000000000000010001000000000000000100000000000000000000000000010000000000010000000000000000,
		120'b00000000000000000000000100000001000000000000000000010000000000000000000100000001000000000000000000000000,
		120'b00000000000000000000000100010010000100000000000000000000000100000000000000000000000000010000000000000000,
		120'b00000000000000000000000000000000000000000000000100000000000000000000000100000000001000010000000100000000,
		120'b00000000000000000000000100010000000000000000000100010000000000000000000100000000000000010001000100000001,
		120'b00000000000000000000000000010000000000000000000100100000000100000000000100000000000000000000000000000010,
		120'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000001,
		120'b00000000000000000000000000000001000000000000000000010000000000000000000100000001000000010001000000000000,
		120'b00000000000000000000000000010000000000000000000000000000000000010000000000000000000000010000000000000001,
		120'b00000000000000000000000000010001000000000001000100000000000000000000000000000000000000010001000000000000,
		120'b00000000000000000000000000100000000100000000000000100000000000000000000100000000000000100000000000000000,
		120'b00000000000000000000000000000010000100000000000000000000000000000000000000000000000000010010000000000001,
		120'b00000001000000000000000100010000000000000000000100010010000000000000000100000000000000000000000100000000,
		120'b00000000000000010000000000010000000000000000000000010000000000000000001000010000000000000000000000000000,
		120'b00000000000000000000000000100010000000000000000000000000000000000000000000000000000000010000000000000001,
		120'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000010,
		120'b00000000000000010000000000010000000000000000000000010000000000000000000000000000000000000000000000000001,
		120'b00000000000000000000000000000000000000000001000100010000000000000000000000010000000000010000000000000000,
		120'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000010000000000000,
		120'b00000000000000000000000000000001000000000010000000010000000000000000001000010001000000000000000000000000,
		120'b00000000000000000001000000000001001000000000000000000000000000000000000000000000000000110001000000000000,
		120'b00000000000000000000000100010001000000000000000000000000000000000001000000000000000000010000000100010000,
		120'b00000000000000010000000000010000000000000000000000010000000000000000000000000000000000110000000000010000,
		120'b00000000000000000000000100000000000100000000000100000001000000000000000000000000000100000000000000000000,
		120'b00000001000000000000000000000000000000000000000000000001000100000000000100000000000100000000000000000001,
		120'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000100010000000100000000000000000001000000000000000000000000,
		120'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000010001000000010001,
		120'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000010001000100000000,
		120'b00000000000000010000000000000001000000000000000100000000000000000000000000010000000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000,
		120'b00000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000100010001,
		120'b00000000000000000000000000000000000000000000000000000000000000010000000000010000000000010000001000000000,
		120'b00000000000000000000000000000001000000000001000000000000000100000000000100000000000000010000000100000001,
		120'b00000000000000000000000000000001000100000001000000000000000000000000000100000000000000010000000100000000,
		120'b00000000000000010000000000010001000000000000000000000000000000000000000100000000000000100000000000010000,
		120'b00000000000100000000000000000000000000000000000000010000000000000000000100000000000000010001000000000000,
		120'b00000000000000000000000000000000000000000000000000010000000000000000000100000001000000010000000000010000,
		120'b00000000000000010000000000000000000000000000000100010001000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000100000000000000000000000000000001000000000000000000010000000000000000000100000000,
		120'b00000000000000000000000000000001000000000000000000010000000000000000000100000001000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000000000000000100000000000100000000000100010000000000000000,
		120'b00000000000000000000000000000000000000000000000000010000000100010000000100000000000000000000000000000000,
		120'b00000000000000000000000000000000000000000001000100010000000000000000000000000000000000010000000000000000,
		120'b00000001000000000000000000010000000000000000000100000000000000000000000000000000000000000001000000000001,
		120'b00000001000000000000000000010000000000000000001000010000000100000000000000010001000000010000000100000000,
		120'b00000000000000000000000100010001000000000000000100000000000000000000000000010000000000000000000000000000,
		120'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000010000000100000001,
		120'b00000000000000000000000000010000000100000001000100000000000000000001000000000000000000010000000100000000,
		120'b00000000000000000000000000000001000000000000000000000001000000000000000000000000000000010000000000000001,
		120'b00000000000000000000000000000001000000000001000000000000000000000000000000000001000000010000000000000001,
		120'b00000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000,
		120'b00000000000000000001000000000001000100000000000100010000000000000000000100000000000000010000000000000000,
		120'b00000000000000000000000000010001000000000000000100010000000000000000000100000000000000010000000100000000,
		120'b00000000000000010000000000000000000000000000000100010000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000100000000000000000000000100010000000000000000000000000000000100000001000000000000,
		120'b00000000000000000000000000010010000100000001000100000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000100000001000000000000000100000000000000000000000000010000000000010000000000000000,
		120'b00000000000000000000000000010000000100000000000000000000000100000000000000000000000000100001000000000001,
		120'b00000001000000000000000100010001000100000000000000000000000000000000000100000000000000010000000100000000,
		120'b00000000000000000000000000010000000000000000000100000000000000000000000000010000000000000000000000010000,
		120'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000,
		120'b00000001000000000000000100010000000000000000000100010000000000000000000000000000000000000000000100000000,
		120'b00000000000000000000000000000000000100000000000000010001000000000000000100000000000000010000000100000010,
		120'b00000000000000000000000000010000000000000001001000000000000000000000000000010000000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000000000001000000000000000000000001000000010000000000000001,
		120'b00000000000000000000000000000001000100000000000000000010000000000000000000000000000000100000000000010000,
		120'b00000000000000010000000000000000000100000001000100000000000000000000000000000000000000010000000000000000,
		120'b00000000000000010000000000000000000000000000000000000000000100000000000100010000000000010000000000000000,
		120'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000100000001,
		120'b00000000000000010000000000010000000100000000000100010000000000010000000000000000000000010000000000000000,
		120'b00000000000000010000000000000000000000000000000100010000000000000000000000000000000000000001000000000000,
		120'b00000000000000000000000100010000000100000001000100000001000000000000000000000000000000010000000100000000,
		120'b00000001000000000000000000010011000000000000000000000001000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000000010000000100000000000000000000000000000000000000010000000000100000000000000000,
		120'b00000000000000000000000000100000000000000000000100000000000100000000000000000000000000000000000000000001,
		120'b00000000000000000000000000000000000000000001000000000000000100000000000000000000000000010000000100000001,
		120'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000010001000000000000,
		120'b00000000000000010000000000000000000000000000001000010000001000000000000100000001000100000000000000000000,
		120'b00000000000000010000000000000000000000000000001000010000000100000000000000000000000000000010000000000001,
		120'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000000000001000000000000000100010000000000000000000000000000,
		120'b00000000000000010000000100100000000000000000000100000000000000000000000100010000000000000000000000000000,
		120'b00000000000000000000000000000000000100000001000000000000000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000001000000001,
		120'b00000000000000000000000000010000000000000000000000010000000000010000000100010000000000000000000000000000,
		120'b00000000000000000000000000010000000100000000000100010000000000000000000000010000000000000000000000000000,
		120'b00000000000000000000000100000010001000000000000100000000000000000000000000000000000000100000000100000000,
		120'b00000000000000000000000100010000001000000000000000010000000000000000000000000000000000010000000100000000,
		120'b00000000000000000000000000010010000000000001000100000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000000000000000000000000000100000001000000000000000000010000,
		120'b00000000000000000000000000000000000000000000000000000001000000000000000100000000000000010001000000000001,
		120'b00000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000001,
		120'b00000000000000000000000000010000000100000000001000010000000100000000000000000000000000000000000100000000,
		120'b00000000000000010000000000010000000100000000000000000000000000000000000000000000000000010000000000000001,
		120'b00000001000000000000000000010001000100000000000100000000000000000000000100010000000000000000000000000000,
		120'b00000000000000000000000100010001000100000001000000000000000000000000000100000000000000010000000100000000,
		120'b00010000000000000000000000000001000000000000000000000000000000000000000100000000000000010000000000000000,
		120'b00000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000001,
		120'b00000000000000000000000000000001000100000001000100010000000100000000000000000000000000010000000000000001,
		120'b00000000000000000000000000000001000000000000000000010000000000000000000100000000000000010000000100000000,
		120'b00000000000000000000000100000000000000000000000000100000000100000000001000000001000000000001000100000000,
		120'b00000000000000000000000100000000000000000000000000000000000000000000000100000001000000010001000000000000,
		120'b00000000000000000000000000000001000000000001000100000000000000000000000000010000000000000000000000000000,
		120'b00000001000000000000000000010000001000000000000100000000000000000000000100000000000000010001000100000000,
		120'b00000000000000000000000000000000000100000000000100000000000000000000000000000000000000000001000000010001,
		120'b00000000000000000000000000010000000000000000001000010000000100000000000100000000000000000000000100000001,
		120'b00000000000000000000000000000000000000000000000000010000000000000000000000010001000000010000000100000001,
		120'b00000000000000010000000000010000000000000000000000000000000000000000000100010000000000010000000000000000,
		120'b00000000000100000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000000000001000000000000000000000001001000000000000000000000000000000000000000000001,
		120'b00000000000000000000000000010000000100000000000000010000000000000000000100000001000000000000000000000001,
		120'b00000000000000000000000000010000000100000000000000000000000000000000000000000000000000010000000000000001,
		120'b00000000000000000001000000010000000100000000000100100001000000000000000000000001000000100000000000000000,
		120'b00000000000000000000000000000000000100000000000000010000000100000000000100010000000000010001000100000000,
		120'b00000000000000000000000100000000000100000000000000010000000000000000000100000001000000000001000000000000,
		120'b00000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000001,
		120'b00000000000000000000000100010000001000000000000000010000000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000100100010000000000000000000010000000000000000000000000000000000010001000000000000,
		120'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000000001000000000010000100010000000000000000000100010001000000000000000000000000,
		120'b00000000000000000000000100010000000000000000000100010000000000000000000000000000000000000000001000000001,
		120'b00000000000000000000000000010001000000000000000000000001000000000000000100000000000000010000000000000000,
		120'b00000000000000000000000000010010000000000000000000000000000000000000000100000000000000010000000000000000,
		120'b00000000000000000001000000000000000000000000000000000000001000000000000000000000000000100000000000000000,
		120'b00000000000000000000000000010000000000000000000000000000000100000000001000000001000000000001000000000001,
		120'b00000000000000000000000000000000000100000001000100000000000100000000000100000000000100010000000000000000,
		120'b00000000000000000001000100000001000100000001000100000000000000000000000100000000000000010000000000000000,
		120'b00000000000000000000000000000000000100000000000100000001000000000000000000000000000100000000000000000000,
		120'b00000000000000000001000000010001000000000000000000010000000000000000000000000000000000100000000000000000,
		120'b00000000000000000001000000000000000000000000000100000000000100000000000000000000000000010000000000000000,
		120'b00000000000000000000000000000000000000000000000100000000000100000000000000000000000000000001000000000000,
		120'b00000000000000000000000000000000000000000000000100010000000000000001000000010000000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000000010001000000000000000100000000000000000000000000000001,
		120'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000001,
		120'b00000000000000000000000100000001000100000000000100000000000000000000000000010000000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000000000001000000000000000100000001000000010000000000000001,
		120'b00000000000000000000000000100000000100000001000000010001000000000000000000000000000000100001000000000001,
		120'b00000000000000000000000000100000000000000000000000000000000100000000000100000000000000010000000000000000,
		120'b00000000000000000000000000010001000100000001000100010000000000000000001000000000000000010001000100000000,
		120'b00000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000,
		120'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000100000001000100000000000000100000000000000000000100000000000000010000000100000001,
		120'b00000000000000000000000000010000000100000000000100010000000000000000000000010000000000010000000000000001,
		120'b00000001000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000,
		120'b00000000000000000000000000000001000000000000000000000000001000000000000000010000000000000000000000000001,
		120'b00000001000000000000000000010000001000000010000100000000000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000100000001,
		120'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000,
		120'b00000000000000000000000000010001000000000000000000000000001000000000000100000000000000000000000000000000,
		120'b00000001000000000000000000000000000000000000000100010001000000000000000000000000000000010000000000000000,
		120'b00000001000000000000000100010000000000010000000000000000000100000000000100000000000000000000000000000001,
		120'b00000001000000000001000000000000000100000000000000000000000000000000000000000000000000100000000000000000,
		120'b00000000000000000000000000010001000000000000000000010000000100000000001000000001000000000000000000000000,
		120'b00000000000000000000000000100000000000000000000100100000000000000000000000000000000000010000000100000000,
		120'b00000001000000000000000100010000000100000000000100010000000000000000000000000000000000000000000100000000,
		120'b00000000000000000001000000010000000100000001000000000000000000000000000100000000000000010000000000000001,
		120'b00000000000000000000000000100000000000000000000000000000001000000000000100000000000000010000000000000000,
		120'b00000000000000000001000000010001000000000000000000000000000000000000001000000000000000000000000000000000,
		120'b00000000000000000001000000000001000000000000000000000000000000000000000000000000000000010000000000000001,
		120'b00000000000000000000000000010001000000000000001000000000000100000000000000000000000000000000000000000000,
		120'b00000000000000010000000000000000000000000000000100000000000100000000000000000000000000000000000000000000,
		120'b00000001000000000000000000000000000100000001000000000000000100000000000000000000000000010000000000000000,
		120'b00000000000000000000000100010001000100000000000100000001000000000000000000000000000000010000000100000000,
		120'b00000000000000000000000000000000000100000000000000000001000000000000000000000000000000110001000100010000,
		120'b00000000000000000000000000000000000100000001000100000001000000000000000000000000000000010000000100000001,
		120'b00000000000000000001000000000001000000000000000100000001000000000000000100000000000000010000000000000000,
		120'b00000000000000000000000100000000000000000000000000010000000100000000000100000000000000010001000100000000,
		120'b00000000000000000000000000000000000000000000000100000000001000000000000000000001000000100000000100000000,
		120'b00000000000000000001000100000000000000000000000000000000000100000000000000000000000000010000000000000001,
		120'b00000000000000000000000000010000000100000000000000000000000100000000000100000000000000010000000100000001,
		120'b00000001000000000000000000000000000100000000000100000000000000010000000000000000000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000001,
		120'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000100000001,
		120'b00000000000000000000000000000001000000000000000100000000000000000001000000000000000000000000000000010000,
		120'b00000000000000000001000000000000000100000001000100000000000000000000000100000000000000010001000000000000,
		120'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000,
		120'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000100000001000000000000,
		120'b00000000000000000000000100000001000100000000000100000000000000000000000000000000000000010000000100000000,
		120'b00000000000000000000000100010000000100000000000100000000000000000000000000010000000000000000000000000001,
		120'b00000000000000000000000000010000000100000000000000010000000000000000000100000000001000100001000000000000,
		120'b00000000000000000000000000000010000100000001000000000000000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000000000000100000000000000010000000100000000000000000000000000010000000000000001,
		120'b00000000000000000000000000000001000000000000000000000000000100000000000000000000000000010000000000000001,
		120'b00000000000000000000000100000000000100000000000100010000000000000000000000000000000000000001000000000001,
		120'b00000000000000000000000000010000000100000001000000010000000000000000000100000000000000000000000000000000,
		120'b00000000000000000000000100000001000100000000000100000000000000000000000000000000000000010000000100000000,
		120'b00000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000010000,
		120'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000100000011,
		120'b00000000000000000000000000000010000100000001000100000000000000000000000000000000000000010000000100000000,
		120'b00000000000000000000000000010000000000000000000000010000000000000000000000000000000000100000000000000000,
		120'b00000000000000000000000000000000000100000000001000000001000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000010001000000000000000100000000000000010000000000000000000000000000000100000000,
		120'b00000000000000000000000000010000000100000000000000100000000000000000001000000001000000000000000000000001,
		120'b00000000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000,
		120'b00000000000000000000000000010000000100000000000000000000000000000000000100000000000000010001000100000000,
		120'b00000000000000000000000000010000000000000001000100010000000000000000000100000000000000000000000000000000,
		120'b00000000000000000000000000000000000000000000000100010000000000000001000100000000000000000000000000000000,
		120'b00000000000000000000000000000001000000000000000000010000000000000000000100000000000000100000001000000000,
		120'b00000000000000000000000000000000000000000000000000010001000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000000010001000100000000000100000000000000000000000100000001000000100000000100000001,
		120'b00000000000000000001000000000000000000000000000000010000000000000000000000000000000000010010000100000010,
		120'b00000000000000010000000000010001000000000000000000000000000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000000000010000000000000000000000000000100000000000000000000000000010000000000000001,
		120'b00000000000000000000000000000000000000000000001000000000000100010000000000000000000000000000000000000000,
		120'b00000000000000000000000000000001000000000000000000010000000100000000000100010001000000010000000000000000,
		120'b00000000000000000000000000010000000000000000000000000000000100000000000000000000000100010000000000000000,
		120'b00000000000000000000000000010000000000000000000000000001000000000000000000000000000000010000000000000001,
		120'b00000000000000000000000000100001000000000000000000000000000000000000000000000000000000100000000000000001,
		120'b00000000000100000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000,
		120'b00000000000000000000000000010001000000000000001000100000000000000000001000000000000000000001000100000000,
		120'b00000000000000000000000000010001000000000000000000000000000100000000000000000000000000100000000100000000,
		120'b00000000000000100000000000000001000000000000000100010000000000000000000100000000000000000001000000000000,
		120'b00000000000000000000000000010001000000000001001000000000000000000000000000010000000000000000000000000000,
		120'b00000001000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001,
		120'b00000000000000000000000000010000000100000000000000000000000000000000000000010000000000010001000000000001,
		120'b00000000000000010000000000000000000000000000000000000000000000010000000000000000000000100000000000000000,
		120'b00000001000000000000000000010000000100000000000100000000000000000000000000000001000000010000000100000001,
		120'b00000000000000000000000000010000000000000000000100010000000000000000000000000000000000010000000000000000,
		120'b00000000000000000001000000000000000000000000000000000000000100000000000100000000000000010000000000000000,
		120'b00000000000000000000000000000000000100000000000000000000000100000000000000000001000000010000000000000001,
		120'b00000001000000000000000000000000000100000000000000000000001000000000000000000001000000010000000000000001,
		120'b00000000000000000000000000010000000000000000000000000000000100000000000000000000000000010000000000010001,
		120'b00000000000000000000000000010001001000000000000000000000000000000000000100000001000000100000000000000000,
		120'b00000000000000010001000000000000000100000000000100000000000000000000000000010000000000100000000000000000,
		120'b00000000000000000000000100000000000000000000000000010000000000000001000000000000000000010000000000000000,
		120'b00000000000000000000000000010000000100000000001000000000000000000000000000000000000000010000000100010000,
		120'b00000000000000000001000000000000000100000000000100010001000000000000000000000000000000100000000000010000,
		120'b00000000000000000000000000010000000100000000000000000001000000010000000000000000000000010000000000000001,
		120'b00000001000000000000000000000000001000000000000000000000000100000000000100000000000000000000000000010001,
		120'b00000001000000000000000000000000000100000000000000000000001000000000000000000000000000010000000000000001,
		120'b00000000000000000000000000010000000000000000000100010000000000000000000100000000000000000000000100000001,
		120'b00000000000000000000000000100001000100000000000000000000000000000000000000000000000000000000000000000001,
		120'b00000000000000000000000000000010000100000000000000000000000000000000000100000000000000100000000000000000,
		120'b00000000000000000000000000000000000000000000000100000001000100000000000000000000000000010001000000000000,
		120'b00000000000000000000000100010001000100000000000000000000000000000000000000000000000100100000000000000001,
		120'b00000000000000000000000000000000000100000000000000000000000000000000000100000000000000000000000000000001,
		120'b00000001000000000000000100010001000100000000000000010000000000000000000100000000000000000001000000000000,
		120'b00000000000000000000000000000000000000000001000000010000000100000000000000000000000000000000000000000001,
		120'b00000000000000000000000100000000000000000000000000010001000000000000000000010000000000000000000000000001,
		120'b00000000000000000001000000000000000100000001000100000000000000000000000100000000000000010010000000000000,
		120'b00000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000,
		120'b00000001000000000000000000000001000000000000000000000000000000000000000000000000000000010000000000000000,
		120'b00000000000000000000000100000000001000010000000000000000000000000000000100000000000000100001000000000000,
		120'b00000000000000000000000000000001000000000000000100010000000000000000000000000000000000010001000100000000,
		120'b00000000000000000000000000010000000000000000000100000000000000000000000000010000000000000000000000000000,
		120'b00000000000000000000000000000011000100000000000100000000000000000000000100000000000000100000001000000001,
		120'b00000000000000000000000000010001000000000000000100000000000000000000000000000000000000000000000100000000,
		120'b00000000000000000001000000000000000000000000000100000001000000000000000100000000000000010000000000000000,
		120'b00000000000000000000000100000001000100000000000100000001000000000000000000000000000100000000000000000000,
		120'b00000000000000000000000000000000000100000000000000000001000000000000000000010000000000000000000100000001,
		120'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001,
		120'b00000000000000000000000000010001000100000001000000000001000000000000000000000000000000110000000000010000,
		120'b00000000000000000000000000100000000100000000000000000000000000000000000000000000000000100000000000010000,
		120'b00000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001,
		120'b00000000000000000000000100010010000000010000000100010000000000000000000100000000000000010000000000000000,
		120'b00000001000000000000000100000000000000000000000000000000000100000001000000000000000000000000000000000000,
		120'b00000001000000000000000000000000000000000000001000000000000000000000000000010000000000000000000000000001,
	}
	
	localparam bit [7:0] alphabet [0:25] = '{
		8'b00000010,
		8'b00000011,
		8'b00000100,
		8'b00000101,
		8'b00000110,
		8'b00000111,
		8'b00001000,
		8'b00001001,
		8'b00001010,
		8'b00001011,
		8'b00001100,
		8'b00001101,
		8'b00001110,
		8'b00001111,
		8'b00010000,
		8'b00010001,
		8'b00010010,
		8'b00010011,
		8'b00010100,
		8'b00010101,
		8'b00010110,
		8'b00010111,
		8'b00011000,
		8'b00011001,
		8'b00011010,
		8'b00011011,
	}
	
	// local parameters
	localparam S_IDLE = 0;
	localparam S_CALC = 1;
	localparam S_DONE = 2;
	
	// logics
	logic [1:0] state_r, state_w;
	logic finish_r, finish_w;
	logic [103:0] word_count_r, word_count_w;
	logic [119:0] word_r, word_w;
	logic similarity_word_w        [0:COUNT_DICT_SIZE - 1]
	logic similarity_word_r        [0:COUNT_DICT_SIZE - 1]
	logic [4:0] similarity_value_w [0:COUNT_DICT_SIZE - 1]
	logic [4:0] similarity_value_r [0:COUNT_DICT_SIZE - 1]
	logic [4:0] max_similarity_value_r, max_similarity_value_w;
	
	interger i;
	
	// assign values
	assign o_similarity_finished = finish_r;
	initial begin
		for (i = 0; i < COUNT_DICT_SIZE; i = i + 1) begin
			assign o_similarity_word[i] = similarity_word_r[i];
		end
	end
	
	always_comb begin
		state_w = state_r;
		finish_w = finish_r;
		word_count_w = word_count_r;
		word_w = word_r;
		max_similarity_value_w = max_similarity_value_r;
		
		initial begin
			for (i = 0; i < COUNT_DICT_SIZE; i = i + 1) begin
				similarity_word_w[i] = similarity_word_r[i];
				similarity_value_w[i] = similarity_value_r[i];
			end
		end
		
		case (state_r)
			S_IDLE: begin
				if (i_start) begin
					state_w = S_CALC
				end
			end
			S_CALC: begin
                interger ptr_word;
                interger charac;
                initial begin
                    for (charac = 0; charac < 26; charac = charac + 1) begin
                        initial begin
                            for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
                                if (alphabet == i_word[ptr_word:ptr_word + 7]) begin
                                    word_count_w = word_count_w + charac * 16
                                end
                            end
                        end
                    end
                end

                interger wd;
                initial begin
                    for (wd = 0; wd < COUNT_DICT_SIZE; wd = wd + 1) begin
                        initial begin
                            for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 4) begin
                                // output the smaller value
                                if (count_dict[ptr_word:ptr_word + 3] >= word_count[ptr_word:ptr_word + 3]) begin
                                    similarity_value_w[wd] = similarity_value_w[wd] + word_count[ptr_word:ptr_word + 3]
                                end else begin
                                    similarity_value_w[wd] = similarity_value_w[wd] + count_dict[ptr_word:ptr_word + 3]
                                end
                            end
                            
                            if (similarity_value_w[wd] > max_similarity_value_w) begin
                                max_similarity_value_w = similarity_value_w[wd]
                            end

                        end
                    end
                end

                ptr_word = 0;
                initial begin
                    for (i = max_similarity_value_w; i >= 0; i--) begin
                        if (ptr_word >= 20) begin
                            break
                        end
                        initial begin
                            for (wd = 0; wd < COUNT_DICT_SIZE; wd = wd + 1) begin
                                if (ptr_word >= 20) begin
                                    break
                                end
                                if (similarity_value_w[wd] == max_similarity_value_w) begin
                                    similarity_word_w[ptr_word] = 0'b1
                                    ptr_word = ptr_word + 1
                                end
                            end
                        end
                        max_similarity_value_w = max_similarity_value_w - 1
                    end
                end
                
				state_w = S_DONE;
				finish_w = 1'b1;
			end
			S_DONE: begin
				finish_w = 1'b0;
				state_w = S_IDLE;
			end
		endcase
		
	end

	always_ff @ (posedge i_clk or negedge i_rst_n) begin
		if (!i_rst_n) begin
			finish_r <= 0;
			state_r <= S_IDLE;
			word_count_r <= 104'b0;
			word_r <= 120'b0
			max_similarity_value_r <= 4'b0;
			initial begin
				for (i = 0; i < 500; i = i + 1) begin
					count_dict[i] = 104'b0;
				end
			end
			initial begin
				for (i = 0; i < 26; i = i + 1) begin
					alphabet[i] = 8'b0;
				end
			end
			initial begin
				for (i = 0; i < COUNT_DICT_SIZE; i = i + 1) begin
					similarity_value_r[i] = 1'b0;
					similarity_value_r[i] = 120'b0;
				end
			end
		end else begin
			finish_r <= finish_w;
			state_r <= state_w;
			word_count_r <= word_count_w;
			word_r <= word_w;
			max_similarity_value_r <= max_similarity_value_w;
			initial begin
				for (i = 0; i < COUNT_DICT_SIZE; i = i + 1) begin
					similarity_word_r[i] = similarity_word_w[i];
					similarity_value_r[i] = similarity_value_w[i];
				end
			end
		end
	end
endmodule

module Viterbi (
    input i_clk,
    input i_rst_n,
    input i_start,
    input i_next,
    input [31:0] i_prob[0:2],
    input [4:0] i_char[0:2],
    output [119:0] o_seq,
    output o_stepped,
    output o_finished
);
    localparam S_IDLE = 2'd0;
    localparam S_CALC = 2'd1;
    localparam S_TOP = 2'd2;
    localparam S_DONE = 2'd3;

    localparam [15:0] transition_prob[0:728] = '{
        16'h0235,
        16'h00fa,
        16'h0164,
        16'h00ca,
        16'h009c,
        16'h00f8,
        16'h0074,
        16'h00b6,
        16'h0147,
        16'h0033,
        16'h0024,
        16'h009f,
        16'h00f9,
        16'h0097,
        16'h0136,
        16'h013a,
        16'h0010,
        16'h00c7,
        16'h01aa,
        16'h0270,
        16'h0056,
        16'h003e,
        16'h00e6,
        16'h0009,
        16'h0045,
        16'h0007,
        16'h0000,
        16'h0002,
        16'h0034,
        16'h006f,
        16'h0054,
        16'h0003,
        16'h0010,
        16'h0041,
        16'h0006,
        16'h0049,
        16'h0002,
        16'h0017,
        16'h00ee,
        16'h004f,
        16'h017e,
        16'h0001,
        16'h0031,
        16'h0002,
        16'h0100,
        16'h0095,
        16'h012b,
        16'h0020,
        16'h002b,
        16'h000b,
        16'h0006,
        16'h003c,
        16'h0006,
        16'h00b2,
        16'h0033,
        16'h0003,
        16'h0002,
        16'h0000,
        16'h0061,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0021,
        16'h0004,
        16'h0000,
        16'h0035,
        16'h0003,
        16'h0001,
        16'h0036,
        16'h0000,
        16'h0000,
        16'h001d,
        16'h000e,
        16'h0002,
        16'h002b,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0022,
        16'h0000,
        16'h0018,
        16'h0085,
        16'h0000,
        16'h0013,
        16'h0003,
        16'h008e,
        16'h0000,
        16'h0000,
        16'h0082,
        16'h0038,
        16'h0000,
        16'h0035,
        16'h002c,
        16'h0001,
        16'h0001,
        16'h00bd,
        16'h0001,
        16'h0000,
        16'h0025,
        16'h000c,
        16'h006c,
        16'h0024,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h000e,
        16'h0000,
        16'h0039,
        16'h003e,
        16'h0003,
        16'h0002,
        16'h0010,
        16'h00a8,
        16'h0001,
        16'h0006,
        16'h0001,
        16'h006b,
        16'h0001,
        16'h0000,
        16'h0007,
        16'h0004,
        16'h0002,
        16'h0032,
        16'h0001,
        16'h0000,
        16'h0015,
        16'h0021,
        16'h0001,
        16'h0022,
        16'h000b,
        16'h0003,
        16'h0000,
        16'h0009,
        16'h0000,
        16'h01b3,
        16'h009a,
        16'h0016,
        16'h006e,
        16'h00c5,
        16'h0054,
        16'h001a,
        16'h001f,
        16'h0005,
        16'h0019,
        16'h0000,
        16'h0006,
        16'h007f,
        16'h0055,
        16'h0116,
        16'h0011,
        16'h0026,
        16'h000b,
        16'h01b1,
        16'h0143,
        16'h0067,
        16'h0008,
        16'h0032,
        16'h0032,
        16'h0031,
        16'h0019,
        16'h0001,
        16'h03b1,
        16'h0021,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h002f,
        16'h001e,
        16'h0000,
        16'h0000,
        16'h0046,
        16'h0000,
        16'h0000,
        16'h000e,
        16'h0000,
        16'h0000,
        16'h0072,
        16'h0000,
        16'h0000,
        16'h0032,
        16'h0001,
        16'h0012,
        16'h0015,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0002,
        16'h0000,
        16'h009a,
        16'h0029,
        16'h0001,
        16'h0000,
        16'h0001,
        16'h0069,
        16'h0000,
        16'h0005,
        16'h0029,
        16'h0026,
        16'h0000,
        16'h0000,
        16'h000d,
        16'h0002,
        16'h0010,
        16'h0021,
        16'h0000,
        16'h0000,
        16'h002b,
        16'h000f,
        16'h0004,
        16'h0015,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0007,
        16'h0000,
        16'h00b7,
        16'h008b,
        16'h0001,
        16'h0000,
        16'h0001,
        16'h0175,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0078,
        16'h0000,
        16'h0000,
        16'h0003,
        16'h0002,
        16'h0008,
        16'h0079,
        16'h0001,
        16'h0000,
        16'h000f,
        16'h0003,
        16'h001b,
        16'h000d,
        16'h0000,
        16'h0001,
        16'h0000,
        16'h0009,
        16'h0000,
        16'h0082,
        16'h0047,
        16'h0015,
        16'h00ab,
        16'h0041,
        16'h0060,
        16'h0027,
        16'h003c,
        16'h0000,
        16'h0003,
        16'h0000,
        16'h000a,
        16'h0071,
        16'h0037,
        16'h01f9,
        16'h00b1,
        16'h001f,
        16'h0002,
        16'h003e,
        16'h00ce,
        16'h00de,
        16'h0003,
        16'h003a,
        16'h0000,
        16'h0005,
        16'h0000,
        16'h000d,
        16'h0037,
        16'h000f,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h000e,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0001,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0011,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h000f,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0003,
        16'h0008,
        16'h0001,
        16'h0000,
        16'h0000,
        16'h0034,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h001e,
        16'h0000,
        16'h0000,
        16'h0003,
        16'h0001,
        16'h0007,
        16'h0004,
        16'h0000,
        16'h0000,
        16'h0001,
        16'h0015,
        16'h0001,
        16'h0001,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0002,
        16'h0000,
        16'h004f,
        16'h007a,
        16'h0003,
        16'h0004,
        16'h0029,
        16'h00c5,
        16'h0007,
        16'h0002,
        16'h0000,
        16'h00a4,
        16'h0000,
        16'h0004,
        16'h0084,
        16'h0005,
        16'h0001,
        16'h0065,
        16'h0009,
        16'h0000,
        16'h0002,
        16'h0027,
        16'h001d,
        16'h001f,
        16'h0005,
        16'h0001,
        16'h0000,
        16'h003d,
        16'h0000,
        16'h00e5,
        16'h0091,
        16'h001a,
        16'h0002,
        16'h0001,
        16'h00bf,
        16'h0001,
        16'h0000,
        16'h0000,
        16'h0046,
        16'h0000,
        16'h0000,
        16'h0002,
        16'h001b,
        16'h0001,
        16'h004d,
        16'h0032,
        16'h0000,
        16'h0001,
        16'h0019,
        16'h0001,
        16'h0018,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h000e,
        16'h0000,
        16'h0068,
        16'h005b,
        16'h0002,
        16'h004d,
        16'h00ed,
        16'h00ad,
        16'h0016,
        16'h00d0,
        16'h0002,
        16'h0051,
        16'h0002,
        16'h0013,
        16'h0013,
        16'h0006,
        16'h0017,
        16'h005a,
        16'h0001,
        16'h0000,
        16'h0002,
        16'h006a,
        16'h00e3,
        16'h0017,
        16'h000b,
        16'h0001,
        16'h0000,
        16'h0016,
        16'h0001,
        16'h01c7,
        16'h0014,
        16'h0017,
        16'h002a,
        16'h0031,
        16'h0008,
        16'h0093,
        16'h0020,
        16'h0005,
        16'h0011,
        16'h0003,
        16'h0016,
        16'h0056,
        16'h0082,
        16'h0177,
        16'h003d,
        16'h0040,
        16'h0000,
        16'h0139,
        16'h0040,
        16'h0063,
        16'h00bc,
        16'h002a,
        16'h0046,
        16'h0006,
        16'h0009,
        16'h0001,
        16'h00d5,
        16'h005b,
        16'h0000,
        16'h0003,
        16'h0004,
        16'h005f,
        16'h0000,
        16'h0001,
        16'h001c,
        16'h0023,
        16'h0000,
        16'h0000,
        16'h003f,
        16'h000a,
        16'h0000,
        16'h0057,
        16'h0022,
        16'h0000,
        16'h0074,
        16'h0010,
        16'h0016,
        16'h001a,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0007,
        16'h0000,
        16'h003f,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0020,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0004,
        16'h00a0,
        16'h0006,
        16'h0028,
        16'h002f,
        16'h018f,
        16'h0007,
        16'h0015,
        16'h0002,
        16'h00ae,
        16'h0000,
        16'h001b,
        16'h0013,
        16'h0028,
        16'h0027,
        16'h00a5,
        16'h0009,
        16'h0000,
        16'h0018,
        16'h0063,
        16'h005d,
        16'h001e,
        16'h0017,
        16'h0003,
        16'h0000,
        16'h003a,
        16'h0000,
        16'h0166,
        16'h0035,
        16'h0004,
        16'h0029,
        16'h0004,
        16'h00d1,
        16'h0003,
        16'h0001,
        16'h0045,
        16'h0081,
        16'h0000,
        16'h000c,
        16'h000d,
        16'h000c,
        16'h0003,
        16'h0052,
        16'h002c,
        16'h0002,
        16'h0002,
        16'h005c,
        16'h00fe,
        16'h0040,
        16'h0001,
        16'h0008,
        16'h0000,
        16'h000e,
        16'h0000,
        16'h0309,
        16'h0085,
        16'h0002,
        16'h000a,
        16'h0002,
        16'h012c,
        16'h0002,
        16'h0001,
        16'h01c5,
        16'h011d,
        16'h0000,
        16'h0000,
        16'h0011,
        16'h0009,
        16'h0003,
        16'h00de,
        16'h0002,
        16'h0000,
        16'h005f,
        16'h005b,
        16'h0023,
        16'h0035,
        16'h0002,
        16'h0010,
        16'h0000,
        16'h0033,
        16'h0001,
        16'h01e1,
        16'h001c,
        16'h0019,
        16'h0025,
        16'h0016,
        16'h0020,
        16'h0004,
        16'h0014,
        16'h0000,
        16'h001a,
        16'h0000,
        16'h0003,
        16'h003a,
        16'h0024,
        16'h0056,
        16'h0003,
        16'h0022,
        16'h0000,
        16'h0085,
        16'h0071,
        16'h0052,
        16'h0000,
        16'h0001,
        16'h0000,
        16'h0002,
        16'h0006,
        16'h0001,
        16'h0026,
        16'h0025,
        16'h0000,
        16'h0000,
        16'h0003,
        16'h009d,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0058,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h000d,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0001,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0009,
        16'h003a,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0044,
        16'h0000,
        16'h0000,
        16'h002b,
        16'h004b,
        16'h0000,
        16'h0000,
        16'h0002,
        16'h0000,
        16'h0010,
        16'h0029,
        16'h0000,
        16'h0000,
        16'h0006,
        16'h0015,
        16'h0001,
        16'h0000,
        16'h0000,
        16'h0002,
        16'h0000,
        16'h0001,
        16'h0000,
        16'h003f,
        16'h0005,
        16'h0000,
        16'h0005,
        16'h0000,
        16'h0005,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0006,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h000b,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h000c,
        16'h0001,
        16'h0000,
        16'h0000,
        16'h0001,
        16'h0001,
        16'h0000,
        16'h001c,
        16'h0006,
        16'h0002,
        16'h0003,
        16'h0002,
        16'h0015,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0005,
        16'h0000,
        16'h0000,
        16'h0005,
        16'h0006,
        16'h0004,
        16'h0037,
        16'h0007,
        16'h0000,
        16'h0006,
        16'h0018,
        16'h0004,
        16'h0000,
        16'h0000,
        16'h0002,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0149,
        16'h0005,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h000b,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0005,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0003,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0001,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0000,
        16'h0001,
        16'h0006,
    };

    logic [4:0] prev_char_r[0:2], prev_char_w[0:2];
    logic [1:0] state_r, state_w;
    logic [31:0] topN_prob0_r, topN_prob0_w, topN_prob1_r, topN_prob1_w, topN_prob2_r, topN_prob2_w;
    logic [31:0] tmp_prob0_r, tmp_prob0_w, tmp_prob1_r, tmp_prob1_w, tmp_prob2_r, tmp_prob2_w;
    logic [31:0] this_prob_r[0:2], this_prob_w[0:2];
    logic [119:0] tmp_seq_r[0:2], tmp_seq_w[0:2];
    logic [119:0] topN_seq0_r, topN_seq0_w, topN_seq1_r, topN_seq1_w, topN_seq2_r, topN_seq2_w;
    logic [119:0] top_seq_r, top_seq_w;
    logic [4:0] counter_r, counter_w;
    logic stepped_r, stepped_w, finish_r, finish_w;

    assign o_prob[0] = topN_prob0_r;
    assign o_prob[1] = topN_prob1_r;
    assign o_prob[2] = topN_prob2_r;
    assign o_seq = top_seq_r;

    assign o_stepped = stepped_r;
    assign o_finished = finish_r;

    always_comb begin
        state_w = state_r;
        topN_prob0_w = topN_prob0_r;
        topN_prob1_w = topN_prob1_r;
        topN_prob2_w = topN_prob2_r;
        topN_seq0_w = topN_seq0_r;
        topN_seq1_w = topN_seq1_r;
        topN_seq2_w = topN_seq2_r;
        top_seq_w = top_seq_r;

        case (state_r)
            S_IDLE: begin
                if (i_start) begin
                    state_w = S_CALC;
                    topN_prob0_w = 32'b0;
                    topN_prob1_w = 32'b0;
                    topN_prob2_w = 32'b0;
                    topN_seq0_w = 90'b0;
                    topN_seq1_w = 90'b0;
                    topN_seq2_w = 90'b0;
                end
                if (i_next) begin
                    state_w = S_CALC;
                end
                counter_w = 0;
            end
            S_CALC: begin
                if (topN_seq0_r == 0) begin
                    topN_prob0_w = i_prob[0] * transition_prob[i_char[0]];
                    topN_prob1_w = i_prob[1] * transition_prob[i_char[1]];
                    topN_prob2_w = i_prob[2] * transition_prob[i_char[2]];
                    topN_seq0_w = {112'b0, i_char[0]};
                    topN_seq1_w = {112'b0, i_char[1]};
                    topN_seq2_w = {112'b0, i_char[2]};
                    state_w = S_REST;
                    prev_char_w = i_char;
                end else begin
                    if (counter_r < 4) begin
                        if (counter_r < 3) begin
                            tmp_prob0_w = topN_prob0_r * i_prob[counter_w] * transition_prob[(prev_char_r[0] + 1) * 27 + i_char[counter_r]];
                            tmp_prob1_w = topN_prob1_r * i_prob[counter_w] * transition_prob[(prev_char_r[1] + 1) * 27 + i_char[counter_r]];
                            tmp_prob2_w = topN_prob2_r * i_prob[counter_w] * transition_prob[(prev_char_r[2] + 1) * 27 + i_char[counter_r]];
                        end
                        if (counter_r > 0) begin
                            if (tmp_prob0_r > tmp_prob1_r & tmp_prob0_r > tmp_prob2_r) begin
                                tmp_seq_w[counter_r]   = {topN_seq0_r[111:0], 3'b0, i_char[counter_r] + 1};
                                this_prob_w[counter_r] = tmp_prob0_w;
                            end else if (tmp_prob1_r > tmp_prob0_r & tmp_prob1_r > tmp_prob2_r) begin
                                tmp_seq_w[counter_r]   = {topN_seq1_r[111:0], 3'b0, i_char[counter_r] + 1};;
                                this_prob_w[counter_r] = tmp_prob1_w;
                            end else if (tmp_prob2_r > tmp_prob0_r & tmp_prob2_r > tmp_prob1_r) begin
                                tmp_seq_w[counter_r]   = {topN_seq2_r[111:0], 3'b0, i_char[counter_r] + 1};;
                                this_prob_w[counter_r] = tmp_prob2_w;
                            end
                        end
                        counter_w = counter_r + 1;
                    end else begin
                        topN_prob0_w = this_prob_r[0];
                        topN_prob1_w = this_prob_r[1];
                        topN_prob2_w = this_prob_r[2];
                        topN_seq0_w = tmp_seq_r[0];
                        topN_seq1_w = tmp_seq_r[1];
                        topN_seq2_w = tmp_seq_r[2];
                        state_w = S_TOP;
                        counter_w = 0;
                    end
                end
            end
            S_TOP: begin
                if (topN_prob0_r > topN_prob1_r & topN_prob0_r > topN_prob2_r) begin
                    top_seq_w = topN_seq0_r;
                end else if (topN_prob1_r > topN_prob0_r & topN_prob1_r > topN_prob2_r) begin
                    top_seq_w = topN_seq1_r;
                end else if (topN_prob2_r > topN_prob0_r & topN_prob2_r > topN_prob1_r) begin
                    top_seq_w = topN_seq2_r;
                end
                state_w = S_IDLE;
            end
        endcase
    end

    always_ff @ (posedge i_clk or negedge i_rst_n) begin
        if (!i_rst_n) begin
            prev_char_r <= '{3{5'b0}};
            state_r <= S_IDLE;
            topN_prob0_r <= 32'b0;
            topN_prob1_r <= 32'b0;
            topN_prob2_r <= 32'b0;
            tmp_prob0_r <= 32'b0;
            tmp_prob1_r <= 32'b0;
            tmp_prob2_r <= 32'b0;
            this_prob_r <= '{3{32'b0}};
            tmp_seq_r <= '{3{32'b0}};
            topN_seq0_r <= 120'b0;
            topN_seq1_r <= 120'b0;
            topN_seq2_r <= 120'b0;
            top_seq_r <= 120'b0;
            counter_r <= 5'b0;
            stepped_r <= 1'b0;
            finish_r <= 1'b0;
        end 
        else begin
            prev_char_r <= prev_char_w;
            state_r <= state_w;
            topN_prob0_r <= topN_prob0_w;
            topN_prob1_r <= topN_prob1_w;
            topN_prob2_r <= topN_prob2_w;
            tmp_prob0_r <= tmp_prob0_w;
            tmp_prob1_r <= tmp_prob1_w;
            tmp_prob2_r <= tmp_prob2_w;
            this_prob_r <= this_prob_w;
            tmp_seq_r <= tmp_seq_w;
            topN_seq0_r <= topN_seq0_w;
            topN_seq1_r <= topN_seq1_w;
            topN_seq2_r <= topN_seq2_w;
            top_seq_r <= top_seq_w;
            counter_r <= counter_w;
            stepped_r <= stepped_w;
            finish_r <= finish_w;
        end       
    end

endmodule

`timescale 1ns / 100ps
module Dictionary(
	input          i_clk,
	input          i_rst_n,
	input          i_start,
	input  [119:0] i_word,
	output         o_finish,
	output [119:0] o_word,
	output [1:0]   o_state
);
	parameter DICT_SIZE = 500;
	localparam bit [119:0] dict [0:DICT_SIZE - 1] = '{
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000100110001000000011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000100100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000111100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110001000000000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101000000100000100100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000010100000100100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000101010000101000011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100001000000011010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010001000000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100001001100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000100000001001100000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011000101100001000000011010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010000110100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000101110000001000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000011000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000100110001000000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000001000011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000011010000101000011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011100001000000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000001000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100010110000100000000001100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000010000000001000010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000001000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000010010000010000010011000000100000011000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001100001001100000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010001011000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110001011000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000111100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000110000010010001010100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001111,
		120'b000000000000000000000000000000000000111100010000000010100001010100000010000011100001001100010000000001110000111100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011100000101000010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010000001100000100100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000101010000101000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100000001000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101000000100000100100011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000100000010100000100100011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100001010000001100000100100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000110000000011000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010001011000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100001010000010110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100000111100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000010011000001100000100100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010000011010000111100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000101000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000001100000100100011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000010101000001000000001000010101000011110001000000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000100110000011000001001,
		120'b000000000000000000000000000000000000000000000000000000000001010000010100000001100000111100001010000101000001011000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000100100011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011000011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000101000000110100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001000000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000011010000011000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000011000001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000001100000101000010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001100000111100001010000011010000111100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100010100000100110000101000000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000001100000011000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001101000101100001000000011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001000000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000100110000011000011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100,
		120'b000000000000000000000000000000000000000000000000000000000001010000000110000001000000101000010111000100110000011000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011100001000000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000010100000001100000100100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000100000010100000110100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001010100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011000000101000001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000110000001000000101000010111000100110000011000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000100000100100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000011110000101000000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000100000010100001001100010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000101010000001000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000001000000001000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000000010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001100000110100010001000100000000011000010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000001000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101000101000000101000001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011100000001000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101000101000001011000001011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011000001100001011100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000010101000000100001010100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011000000100000011000011010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100000001000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000101010000111100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100001010000000100000111000000110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001100000010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000010010001010100001101000000100000011000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001101000100110001000000011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101000110010000011000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001100001010000010110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000100110001000000011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101000101000000001000001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101000101000001000000001110,
		120'b000000000000000000000000000000000000000000000000000000000001010000010101000001000001011000000101000100000001001100010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001010000101000001011000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100001011000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000101010000001000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011000000001000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000001100000100100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010000110100010110000100000000100100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000010101000001000001011000000101000100000001001100010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000011100000011000010101000101000001101000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101000101000001000000010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110000011000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010000101010000101000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000110100000010000001010000011010001000000010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110000011000000011000011100001011000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000001000001011000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001100001010000000010000001100000110100010001,
		120'b000000000000000000000000000000000000000000000000000001100000110100000011000000100000110100001010000000100001011100000010,
		120'b000000000000000000000000000000000000000000000000000101010000100100001000000010100001001100011010000100010001000000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000010101000100110001000000010001000100010001011000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000110000010000000001000010100000101000000011000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000110000101010000011100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101000101000000011000000011,
		120'b000000000000000000000000000000000000000000000000000000000000011000010011000000100001100000010101000001110001000000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000001100000100100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000001000001011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000100000001000000001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000110000001010000101000010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000011010000011000011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000010011000001100000100100011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000001110000111100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000001010100001001000010000000101000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001000000101000001101000000110001011000010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000001100000100000001000000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000010000000101000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000011010001000000010000000010010000010000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000001001000010000001011000010000000100110000100100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000001000000001000000110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000001100000011110000101000001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000100100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000110000000011000001010000101110000011000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010011000000100000011000011010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000110000001010001001100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010000100110000011000010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000011010000001000000001000010111000010100001001100010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000100000001000000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000001110000001100001010100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000011010000011110000001000010001000011100001000000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000100000011000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010110000100000001001100001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010000011000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000001100000011000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010000011110000001000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011000001100001010000010110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000010100000001000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000001100001000000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000011000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000110000001010000111100010110,
		120'b000000000000000000000000000000000000000000000000000000000000000000001101000000100001001100000110000011110000011000001000,
		120'b000000000000000000000000000000000000000000000000000000000000100100000100000100110000001000000110000101000000011000010011,
		120'b000000000000000000000000000000000000000000011010000101010000101000010100000100110000011000010111000010100000111100010110,
		120'b000000000000000000000000000000000000000000000000000000000000000000011010000100110000001000010110000011110000001000001011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000010100000001000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000011010001011000000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000001000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000010100000110000000011000001010000101110000011000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000001110000000100001001100001000000100000001001100010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001110000101000001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000100000000111100001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000110000011100000001000001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100000001000011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000110100000001000000101,
		120'b000000000000000000000000000000000000000000010101000011110000011000001110000001100000100000000010000011110000001000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101000100110000001000010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001101000101100001000000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100000010000001100001001100001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010000011000010101000010100000111100010110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100000110000101010001000000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000000100000011000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000001100001010100001010,
		120'b000000000000000000001101000000100000111100010000000010100001010100000010000011110001001100000110000101010000111100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110000011000010101000011110000011000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010000000100000001100000110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101000101000001011000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000010011000100000001010100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000011010000011000010111000000100001001100010101,
		120'b000000000000000000000000000000000000000000000000000000000001010000010101000011110000011000001110000011100001000000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001010000001000001110,
		120'b000000000000000000000000000000000001010100001111000001100000111000010001000100000000110100000110000101110000011000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000101010001001100010000000100010000011000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000011100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110000011000000011000011100000011000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000010100000011010000101000000010000101010000011000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011110000101000001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000001110000100110000011000010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001100001001100010000000001110000011000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000000110100000110000101010001000000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000101000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000011110000011000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100001001000010000000101000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000100010001101000010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000110000101000001011000000010000001000000011000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100000010000001000001000000001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000010100000100000000100100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001111000010100001010000010110,
		120'b000000000000000000000000000000000000000000000000000000000000000000010100000101010000110100010110000101000000011000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001100000010000001010000001110000011100010000,
		120'b000000000000000000000000000000000000000000000000000011110001000000001010000101010000001000000100000101100000010100000110,
		120'b000000000000000000000000000000000000000000000000000000000000110100000010000011110001000000001010000101010000001000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110000001000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000011110000100000001010000101000000011000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011000000001000010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010000011000010101000101000001000000010001,
		120'b000000000000000000000000000000000000000000000000000000000001010100000110000011110001001100000110000101010000111100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000010100000101000000011000010011000001010000010100000010,
		120'b000000000000000000000000000000000000000000000000000110100001010100001010000011110001011000001110000011100001000000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000011110000101000001001000101010000101000011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000000011000010101000000100001010100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001100001001100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101000011110000001000011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001111000100000000100100010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010001011100000101,
		120'b000000000000000000000000000000000000000000000000000000000000100000001111000010100001000100010001000010100000100100010100,
		120'b000000000000000000000000000000000000000000000000000000000000010100000110000101110001001100000110000101000000011000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000010101000001000000011000001011000000110001011000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000001111000001100000011000011000000101010000011000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000010110000100110001000000000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000110100000110100001010000011100000001000000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000011110001000000001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000110000101000000001000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001010001000000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000100000000100100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000001100001011100000110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000100000000100000110100000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000100000001100000100100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000001101000000100000101000000100000001100001000100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000000011000000100000010100001001100010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000110000101010000101000010100000000110000011000011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001100100000110000001010000111100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001111000010100000011000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000110000011100001000000011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000001000001011000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000010000000101000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011010000101000000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011110000101000001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000001100001000100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000000010000001010001000000010101,
		120'b000000000000000000000000000000000000000000011010000010000001000000001101000100000000111100001001000001000000011000010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100010101000101100001000000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000101000000001000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000010101000001000000011000001011000100000001001100010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011100000001000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000110000010000000001000010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000010110,
		120'b000000000000000000000000000000000000000000000000000000000000000000001111000100000000101000010100000100110000011000010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000001111000100000000101000010101000001000000011000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110001100000010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100001111000101100001000000000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000001010100010011000100000001000100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000010100000101100001000000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000101000001100001010100000010000011010000011000010011,
		120'b000000000000000000000000000000000000000000000000000000000001101000010101000010100001001100010110000001000000011000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000101010001000000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000110100001010100001111000101100001000000000100,
		120'b000000000000000000000000000000000000000000000000000000000000111100000010000001000000101000010011000001100000111000000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010101000100000000100100010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011100000001000001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000010100000100110000011000000011000011100000011000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000110000110000001000000010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001101000010100000100100011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000100110000001000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000001100000100110001000000011000000101010000011000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000110000001000000000101,
		120'b000000000000000000000000000000000000000000000000000000000001001100000110000101010001011000010001000011100001000000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000010100000011100000011000010101000101000001101000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000110000100110000100100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100000010000101010001000000010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000100000000100000110100010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000111100000110,
		120'b000000000000000000000000000000000000000000000000000010000000111100001010000110000001000000001101000011010001000000000111,
		120'b000000000000000000000000000000000000000000000000000000000000010100000010000100000000110100001111000110000001000000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100000101000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000010101000101100001000000001001000101010000101000011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110000011000010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000001010000000110000001000000010000000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001111000010100000100100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100010101000100110001000000001111,
		120'b000000000000000000000000000000000000000000000000000101000000011000000100000100110001011000010000000101000000011000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000010101000011110000011000010011000100110001011000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010101000101000001000000010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000101000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001010000001010000011000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000001000001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000001101000100000001001100010101000011110001000000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100000110000101010000001000011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000011010000100110001000000010101000101000000101000001001,
		120'b000000000000000000000000000000000000000000000000000000000001010000000110000100110001011000010101000001000000101000010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000110110000101000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010001001100000010,
		120'b000000000000000000000000000000000000000000000000000000000000110100000010000011110001000000010100000100110000011000010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000100000011110000101000010100,
		120'b000000000000000000000000000000000000000000000000000010000000111100001010000001010001011000001101000001000000111100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000101000010100001011000001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100000000100100010100,
		120'b000000000000000000000000000000000000000000000000000110100001001100010000000101010000010000000110000100110000101000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100010011000000100001000000000011,
		120'b000000000000000000000000000000000000000000000000000000000000111100010000000010100001010100000010000001000001000000001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001100000100000001111000000100000100100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000010101000010100000100100011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101000110010000011000010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100001101000000100000111000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000111100001010000101010000001000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000101010000001000010011,
		120'b000000000000000000000000000000000000000000010101000011110000011000001110000011110001001100000110000101110001000000001000,
		120'b000000000000000000000000000000000000000000000000000000000000111100000110000100110000010100001101000010100000100100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000010000000111100001010000100110001011000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001010000010110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000011110001001100010110000101010000011000010011,
		120'b000000000000000000000000000000000000000000000000000000000001010000010101000011110000011000000101000101100001010100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111,
		120'b000000000000000000000000000000000000000000000000000000000000100000001111000010100001000100010001000100000000100100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000010101000011110001011000010000000001000000010000000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000110000011100000101000010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000110000101010000101000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100000110000101110000011000001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000001101000000100001010100001010000010000000101000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000110000011010000101000000111000100000001001100010001,
		120'b000000000000000000000000000000000000000000000000000000000001010000010110000100000000101000010111000001100001001100010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000100110001000000000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000001010100001111000001100001011100000110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000101110001000000001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000110100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000010010001000000001011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000010100000001000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000011010000001000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010011000101100001000000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001000000000100000111000001010,
		120'b000000000000000000000000000000000000000000010101000011110000011000001110000101010001001100000010000100010000011000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001101000101010000101000010101,
		120'b000000000000000000000000000000000000111100010000000010100001010100010001000010100001001100000100000101000000011000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110001000000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010,
		120'b000000000000000000000000000000000000000000000000000001100000010000001111000000100001001100010110000101000000111100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000010011000001100000100100010101000100000000111100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100000100100011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100001101000000100000100100010100,
		120'b000000000000000000000000000000000000000000000000000000000001101000010101000100110000011000010001000100000001001100010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000000100000110100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100001101000010100001010100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000000110000011110001000000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000011010000101010000101000001101000000100001011000010010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000010011000001100001011100000110,
		120'b000000000000000000000000000000000000000000000000000000000000000000001000000011110000101000010101000101000000101000001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000010101000011110000011000010101000011110001000000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000011010000100110001010100001111000101100001000000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000110000101010000001000010111000010100001001100010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001100000110100010101000101010000101000001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100001010000101000000101000010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000101110000001000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000001101000100000001000000010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000001000000001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000001101000100010000011000010011,
		120'b000000000000000000000000000000000000000000000000000000000001001100000110000011100001000000010101000101000001011000000100,
		120'b000000000000000000000000000000000000000000000000000000000001001100000110000000110000111000000110000001000000011000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000110000100110000001000010001000011100001000000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000000011000001010000101110001000000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000110000001010001011000001101000001000000111100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000110000010000000011000001101000011010001000000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000010110000011010000001000010111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000110000011010000010000001010000101010001001100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000100110001000000011010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000001000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000100110000001000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000000110001000000001011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000110000001010000101000010111000100000001001100010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000100000001000000000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001100000010000010011000101100001000000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110001000000001001000101010001011000000010,
		120'b000000000000000000000000000000000000000000000000000101010000111100000110000100110000011000000111000001110000101000000101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010100000001100001001100010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100010011000000100000011000001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011010000001000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010000111100010110000100000001001100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100001111000010100001001100010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001100001010000010011000101100001000000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110001000000001011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000100000010100000010000011110000001000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000010100000101000000011000000100000100000001001100010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000001100000011000010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000100000001000000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000100000100000001010100010100,
		120'b000000000000000000000000000000000000000000000000000000000000100000001111000010100000111100001010000000100001001100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000101010000101000000101000001100001001100000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100001111000010100001000000010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000010100001000000001011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000110000001000000111100000110000010100000010000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000011000001110,
		120'b000000000000000000000000000000000000000000010100000001100000101000010011000100000000100000000110000101010000001000000100,
		120'b000000000000000000000000000000000000000000000000000000000000010100000110000001000000111100000010000101110000010100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101000101000000011000011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000110000011010000001000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000100000001000000001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000001001000101000000101000001101000010000000111100000110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101000001110000011000001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000000100000011000010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001100001010100000010000101010001010000000110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010001000000000011,
		120'b000000000000000000000000000000000000000000010100000011110001000000001010000101010000101000000101000011110001000000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000101010000010000000110000011010000011000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000010100000110000001000000000101000011110000101000011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000001000000010101000100000000100100010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100000001000001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010000001000000110000100110000100100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000001100000011000011000,
		120'b000000000000000000000000000000000000000000000000000000000001101000010011000100000000100000000110000101010000001000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000101010001000000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000101110000101000001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001000000100110000001000001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000011010000100110000011000001101000011010000001000001000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001101000000110000001000010101,
		120'b000000000000000000000000000000000000000000000000000000000001001100000110000101010001010000001010000010000000011000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000010011000001100001011100000110000110000001000000001001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000011110001011000001011,
		120'b000000000000000000000000000000000000000000000000000000000000000000010011000001100000001100010000000101010000010000010000,
		120'b000000000000000000000000000000000000000000000000000000000001001100000110000000110000111000000110000101110001000000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000101010000011000001100000100110000001000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000011010000100110000001000010011000000110000101000001101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000110100000110100001101000000100000011000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000011110001000000001010000101010000010000000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100010011000000100001010100010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000000011000001010000100110000011000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100000110000001010001000000001110,
		120'b000000000000000000000000000000000000000000000000000000000001010000000110000100110001011000010101000000100000011000000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110000101000000010,
		120'b000000000000000000000000000000000000000000000000000000000001101000010011000101010001010000010110000001010000111100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000100000110100010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000010000011100001011000001001,
		120'b000000000000000000000000000000000000000000000000000000000000010100000110000001010000101000010111000100000001001100010001,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000000011000011010,
		120'b000000000000000000000000000000000000000000000000000000000000010100000110000100110000101000010110000100100000011000010011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000001010000111100010000000001000000011000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010001000000001001,
		120'b000000000000000000000000000000000001010000000110000010100001001100010000000101000001010000000110000001000000010000000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101000101000001000000000100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001010000101110001000000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000101000000111000010110000100110001000000000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000100000100110000001000001110,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000001101,
		120'b000000000000000000000000000000000000000000000000000100110000011000000011000011100000011000010101000100010000011000010100,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000100110000011000010101000101010000011000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100000001000010100,
		120'b000000000000000000000000000000000000000000000000000101000000111100010000000010100001010100010100000001100001011000010010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010000011010001011000001011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000010010000001000011010
	};
	
	localparam S_IDLE = 2'd0;
	localparam S_CALC = 2'd1;
	localparam S_DONE = 2'd2;
	
	logic [1:0] state_r, state_w;
	logic finish_r, finish_w;
	
	logic similarity_start_r, similarity_start_w;
	wire  similarity_finish_w;
	logic similarity_finish_r, pre_similarity_finish_r;
	wire  [2:0] DTW_state_w; // debug
	logic [2:0] DTW_state_r; // debug
	logic DTW_start_r, DTW_start_w;
	wire  DTW_finish_w;
	logic DTW_finish_r;
	
	wire  similarity_word_w [0:499];
	logic similarity_word_r [0:499];
	logic [119:0] DTW_candidate_word_w [0:19], DTW_candidate_word_r [0:19];
	wire  [119:0] DTW_word_w;
	logic [119:0] DTW_word_r;
	logic [8:0] ptr_r, ptr_w;
	
	integer i;
	assign o_finish = finish_r;
	assign o_word = DTW_word_r;
	assign o_state = state_r;
	
	Similarity sim1(
		.i_similarity_clk(i_clk),
		.i_similarity_rst_n(i_rst_n),
		.i_similarity_start(similarity_start_r),
		.i_similarity_word(i_word),
		.o_similarity_finish(similarity_finish_w),
		.o_similarity_word(similarity_word_w)
	);
	
	DTW dtw1(
		.i_DTW_clk(i_clk),
		.i_DTW_rst_n(i_rst_n),
		.i_DTW_start(DTW_start_r),
		.i_DTW_word(i_word),
		.i_DTW_candidate_word(DTW_candidate_word_r),
		.o_DTW_finish(DTW_finish_w),
		.o_DTW_word(DTW_word_w),
		.o_state(DTW_state_w)
	);
	
	always_comb begin
		state_w = state_r;
		finish_w = finish_r;
		similarity_start_w = similarity_start_r;
		// similarity_finish_w = similarity_finish_r;
		DTW_start_w = DTW_start_r;
		// DTW_finish_w = DTW_finish_r;
		// DTW_word_w = DTW_word_r;
		// DTW_state_w = DTW_state_r;
		DTW_candidate_word_w = DTW_candidate_word_w;
		// similarity_word_w = similarity_word_r;
		ptr_w = ptr_r;
		
		case (state_r)
			S_IDLE: begin
				finish_w = 1'b0;
				if (i_start) begin
					similarity_start_w = i_start;
					state_w = S_CALC;
				end
			end
			S_CALC: begin
				finish_w = DTW_finish_r;
				
				if (similarity_finish_r) begin;
					for (i = 0; i < DICT_SIZE; i = i + 1) begin
						if(similarity_word_r[i] == 1'b1) begin
							DTW_candidate_word_w[ptr_r] = dict[i];
							ptr_w = ptr_r + 1;
						end
					end
				end else if (pre_similarity_finish_r && !similarity_finish_r) begin
					DTW_start_w = 1'b1;
				end
				
				if (finish_r) begin
					state_w = S_DONE;
				end
			end
			S_DONE: begin
				finish_w = 1'b1;
				state_w = S_IDLE;
			end
		endcase
		
	end

	always_ff @ (posedge i_clk or posedge i_rst_n) begin
		if (i_rst_n) begin
			state_r                 <= S_IDLE;
			finish_r                <= 1'b0;
			similarity_start_r      <= 1'b0;
			similarity_finish_r     <= 1'b0;
			pre_similarity_finish_r <= 1'b0;
			DTW_start_r             <= 1'b0;
			DTW_finish_r            <= 1'b0;
			DTW_word_r              <= 120'b0;
			DTW_candidate_word_r    <= '{20{120'b0}};
			DTW_state_r             <= 3'b0; 
			similarity_word_r       <= '{500{1'b0}};
			ptr_r                   <= 9'b0;

			
		end else begin
			state_r                 <= state_w;
			finish_r                <= finish_w;
			similarity_start_r      <= similarity_start_w;
			similarity_finish_r     <= similarity_finish_w;
			pre_similarity_finish_r <= similarity_finish_r;
			DTW_start_r             <= DTW_start_w;
			DTW_finish_r            <= DTW_finish_w;
			DTW_word_r              <= DTW_word_w;
			DTW_candidate_word_r    <= DTW_candidate_word_w;
			DTW_state_r             <= DTW_state_w;
			similarity_word_r       <= similarity_word_w;
			ptr_r                   <= ptr_w;
		end
	end
endmodule

`timescale 1ns / 100ps
module Similarity(
	input          i_similarity_clk,
	input          i_similarity_rst_n,
	input          i_similarity_start,
	input [119:0]  i_similarity_word,
	output         o_similarity_finish,
	output         o_similarity_word [0:499]
);

	parameter COUNT_DICT_SIZE = 500;
	parameter COUNT_SIZE = 26 * 4;

	localparam bit [COUNT_SIZE - 1:0] count_dict [0:COUNT_DICT_SIZE - 1] = '{
		104'b00000000000000010000000000000000000100000000000100000000000000000000000000000000000000000001000000000000,
		104'b00000000000000000000000000010000000000000000000000000000000000000000000000010000000000010000000000000000,
		104'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000100000000000000000000,
		104'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000001,
		104'b00000000000000000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001,
		104'b00000000000000000000000000000000000000000000000000010000000000000000000100000000000000000000000000000000,
		104'b00000000000000000000000000000000000100000000000100000000000000000000000000000000000100000000000000000000,
		104'b00000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000000001,
		104'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000,
		104'b00000000000000000000000000010001000000000000000000000000000000000000000100010000000000000000000000000000,
		104'b00000000000000010000000000010000000000000000000000000000000000000000000100010000000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000,
		104'b00000001000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000,
		104'b00000000000000000000000000010000000000000000000100010000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000,
		104'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000001,
		104'b00000000000000000000000000000000000100000000000100000001000000000000000000000000000100000000000000000000,
		104'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000001,
		104'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001,
		104'b00000001000000000000000100000000000100000000000100000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001,
		104'b00000000000000000001000000000000000000000000000000000000000000000000000000010000000000010000000000000001,
		104'b00000000000000010000000000000000000000000000000000010000000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000000000000000100000000000100000001000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001,
		104'b00000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000001,
		104'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000,
		104'b00000000000000010000000000000000000000000000000000000000001000000000000100000000000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000100000001000000000000000000010000000000010000000000000000,
		104'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000001,
		104'b00000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000100010000000000000000000100000000000000000000000000000000000000000000000000010001,
		104'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000100000000000000000000,
		104'b00000000000000000000000000000000000000000001000000000000000000000000000000000001000000010000000000000001,
		104'b00000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000001,
		104'b00000000000000000000000000000001000100000000000000000000000000000000000000010000000000010000000100000001,
		104'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000100100000000000000000,
		104'b00000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000010000,
		104'b00000000000000000000000100000000000100000000000100000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000100010000000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000000010000000100000000000100000000000000000000000000010000000000010000000000000000,
		104'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001000000000000,
		104'b00000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000010000000100000000001000100001000000000000001000000000000100000000000000000001,
		104'b00000000000000000000000000010000000000000000000000000001000000000000000100000000000000010000000000000000,
		104'b00000001000000000000000000010000000000000000000000000000000000000000000000010000000000010000000000000000,
		104'b00000000000000000000000000010001000000000000000000000000000000000000000100000000000000010000000000000000,
		104'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000,
		104'b00000000000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000,
		104'b00000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001,
		104'b00000000000000010000000000010000000000000000000000000000000000000000000000010000000000000000000000000001,
		104'b00000000000000010000000000000000000000000000000000000000000000000000000100100000000000000000000100000000,
		104'b00000000000000000000000000010000000100000000000000000000000000000000000100010000000000010000000000000000,
		104'b00000000000000010000000000000001000000000000000000010000000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000100010000000000000000000100000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000100000001000000000000000000000000000000000000000000000000000000010000000000000000,
		104'b00000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001,
		104'b00000000000000000000000000010000000100000000000000000000000000000000000000010000000000100000000000000000,
		104'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000100000000000000000,
		104'b00000001000000000000000000000000000000000000000100010000000100000000000000000000000000000000000000000000,
		104'b00000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000000001000000000000000000000000000000000000000100010000000000000000000000000000,
		104'b00000000000000010000000000000000000000000000000000010000000000000000000000010000000000010000000000000000,
		104'b00000000000000000000000000100000000000000000000100010000000000000000000000000000000000000000001000000001,
		104'b00000000000000000000000000000000000100000000000000000000000000000000000000010000000000100000000000000000,
		104'b00000000000000000000000100000011000000000000000000010000000000000000000100000000000000010000000000010000,
		104'b00000000000000010000000000000000000000000000000100000000000000000000000000010000000000000000000000000000,
		104'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000010000,
		104'b00000000000000000000000000000001000000000000000100000000000100000000000000000000000000000000000000000001,
		104'b00000000000000010000000000000000000000000000000100010000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000000000000000000001000000000000000100000000000000010000000000010000000000000000,
		104'b00000000000000000000000000010000000000000000000000000000000000000000000000000001000000010000000000000000,
		104'b00000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000000000,
		104'b00000000000000010001000000000000000000000000000000000000000000000000000100000000000000010000000000000000,
		104'b00000000000000000000000000000000000000000000000100100000000100000000000100000000000000010000000000000000,
		104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000,
		104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000000010001000100000000000000000000000000000000000100000000000100000000000000000000,
		104'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001,
		104'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000100000000000010000,
		104'b00000000000000010000000100000000000000000000000100000000000100000000000000000000000000000001000000000000,
		104'b00000000000000010000000000000000000000000000000100000000000000000000000000010000000000000000000000000000,
		104'b00000000000000010000000000000000000100000000000000000000000000000000000000000000000000100000000000000000,
		104'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000001000000000010000100000000000000000000000000000000000100000000000000100000000100000000,
		104'b00000000000000000000000000000001000000000000000100000001000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000000010001000000000000000000000000000000000000000000010000000000100000000000000000,
		104'b00000000000000000000000000000000000000000000000000000000000100010000000100000000000000000000001000000000,
		104'b00000000000000000000000000010001000000000000000000000000000000000000000100000000000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000000000000000100010000000100000000000000010000000000000000,
		104'b00000000000000000001000000000001000100000000000000000000000000000000000100000000000000100000000100000000,
		104'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000010000000000000000000000010000000000000000000000010000000000000000000000000001,
		104'b00000000000000000000000000000000000000000000000000010000000000000000000100000000000100000001000000000000,
		104'b00000000000000000000000000000000000100000001000000000000000000000000000100000000000000010000000100000000,
		104'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000010001000000000001,
		104'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001,
		104'b00000000000000000000000000010000000000000001000100000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000000000000000000010000100000000000100000000000000000000000000100000000000000000,
		104'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000001,
		104'b00000000000000000000000000010001000000000000000000000000000100000000000100000000000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000000010001000000000000000000000000000000010000000000000001,
		104'b00000000000000000000000100010001000000000000000000000000000000000001000000000000000000000000000000000000,
		104'b00000000000000000001000000000000000100000000000100000000000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000000100001000000000000000000000000000000000000000000000000000000010000000000000001,
		104'b00000001000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000001,
		104'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001,
		104'b00000000000000000000000000010000000000000000000100010000000000000000000100000000000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000000000001000100000000000100000000000000010000000000000001,
		104'b00000000000000010000000000010000000000000000000100000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000010000000000000000000000000000000100000000000000100000000000010000000000000001,
		104'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000,
		104'b00000000000000010000000000000000000100000000000100000000000100000000000000000000000000000001000000000000,
		104'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000,
		104'b00000000000100000000000000010000000000000000000000010000000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000100000001000000000000000000000000000000000000000000000000000000010001000000000000,
		104'b00000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000,
		104'b00000000000000010000000000000000000100000000000100000000000000010000000000000000000000000000000000000000,
		104'b00000000000000000000000000010001000000000000000000000000000100000000000000000000000000000000000000000001,
		104'b00000000000000000000000000010001000000000000000100000001000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000100010001000100000001000100000000000000000000000000000000000000000001000100000000,
		104'b00000000000000000000000100000001000000000000000000000001000000000000000100000000000000000000000100000000,
		104'b00000001000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000010000,
		104'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000010,
		104'b00000000000000000000000000000000000000000000000000000001000000010000000000000000000000010000000000000001,
		104'b00000000000000000000000000010000000000000000000000000001000000000000000000010000000000010000000000000000,
		104'b00000000000000000000000100000001000000000000000100000000000100000000000000010000000000000001000000000000,
		104'b00000000000000000000000100010000000100000001000100000000000000000000000000000000000000000001000100000000,
		104'b00000001000000000000000000010010000000000000000000000001000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000000010001000000000001000100000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000000000000100000000000000000000000000000000000000010000000000010000000000000000,
		104'b00000001000000000000000000010000000000000000000000000000000000000000000100000000000000000000000100000000,
		104'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000001,
		104'b00000001000000000000000000000000000000000001000100000000000100000000000100000000000000000000000100000000,
		104'b00000000000000000000000100000000000100000000000000010001000000000000000000000000000000010000000000010000,
		104'b00000000000000000000000100000001000000000000000000000000000000000000000000010000000000000000000100000000,
		104'b00000000000000000000000000000001000000000001000000000000000100000000000000000000000000100000000000000001,
		104'b00000000000000000001000000000000000000000000000000000000001000000000000100000000000000010000000000010011,
		104'b00000001000000000000000000010000000100000001000100000000000000000000000100010001000000000000000100000000,
		104'b00000000000000000000000100010001000100000010000100000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000000010000000000000000000000001000000000000000000000001000000100000000000000001,
		104'b00000000000000000000000000010000000100000000000000000000000000000000000000000000000100010000000000000001,
		104'b00000000000000000000000000010001000000000000000000000000000000000000000000000000000000010000000000010000,
		104'b00000000000000010000000000010001000100000000000100000000000000000000000000000000000100010000000000000001,
		104'b00000000000000000000000000010000000000000000000000010000000000000000000000010000000000010000000000000000,
		104'b00000000000000000000000000000000000000000000000000010000000000000001000000000000000000000000000000000001,
		104'b00000000000000000000000000000000000000000000001000000000000000000000000000000001000000000001000000000000,
		104'b00000000000000000001000000000000000000000000000100000000000000000000000100000000000000010001000000000000,
		104'b00000000000000010000000000000000000000000000000000000000001000000000000000000000000000010000000000000000,
		104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000,
		104'b00000000000000010000000000000000000100000000000000000000000000000000000000010000000000100000000000000000,
		104'b00000000000000000000000000000000000000000000000100010000000000000000000100000000000100000000000000000000,
		104'b00000000000000000000000000010001000100000000000000000000000000000000000100010001000000000000000000000000,
		104'b00000000000000000000000100000000000000000001000000000000000100000000000100000000000000000000000100010000,
		104'b00000000000000000000000000000001000000000000001000000000000000010000000000000000000000000000000000010000,
		104'b00000000000000000000000000000000000000000000000000000000000000000000000100100001000000000000000000000000,
		104'b00000000000000000000000000000001000000000000001000000000000100000000000000010000000000000000000100000000,
		104'b00000000000000000000000100010000000100000000000100000000000000000000000000100001000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000100000001,
		104'b00000000000000000000000000000001000000000000000000010000000100010000000100000000000000000000000000000000,
		104'b00000000000000000000000000000001000000000000000000000000000000000000000000010000000000010000000000000000,
		104'b00000000000000010001000000000000000100000000000000000000000000000000000100000000000000100000000000000000,
		104'b00000001000000000000000000000001000100000000000000000000000000000000000000000000000000010000000000000001,
		104'b00000000000000000000000000000000001000000000000100000000000000000000000000000000000000010001000000000000,
		104'b00000001000000000001000000000000000100000000000000000000000000000000000000000000000000010000000000000000,
		104'b00000001000000000001000000000000000100000001000000000000000000000000000100000000000000000000000100000001,
		104'b00000000000000000000000000000000000000000000001000000000000000010000000000000000000000000000000000010000,
		104'b00000000000000000000000000010001000000000000000000000001000000000000000100000000000000010000000000000000,
		104'b00000001000000000000000000000000000000000001000100010001000000000000000000000000000000000000000100000001,
		104'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000010001000000000001,
		104'b00000000000000000000000100000000000100000001000100000000000000000000000000000001000000000000000000000000,
		104'b00000000000100000000000000000001000000000000000000000000000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000100001000000000000,
		104'b00000001000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000001,
		104'b00000000000000000000000100000001000100000000000000000000000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000000000001000000000000000000000000000000000000000100000000000000000001000000000001,
		104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000000000,
		104'b00000000000000000000000000000001000000000000000100000000000000000000000000000000000000010001000000000000,
		104'b00000000000000000000000000010001000000000000000000000000000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000100000000000100000000000000010000000000000000000000000000000000010001000000000000,
		104'b00000000000000000000000000000000000100000000000000010000000100000000000000000001000000100000000000000001,
		104'b00000000000000000000000000000001001000000000000000000000000000000000000000010000000000100000000100000001,
		104'b00000001000000000001000100010001000100000000000000010000000000000000001000000000000000010000000000000000,
		104'b00000001000000000000000100000000000100000000000000010000000000000001000000000000000000000000000000000010,
		104'b00000000000000000000000000000000000000000000000000000001000100000000000100000000000000000000000000000001,
		104'b00000000000000000000000100000000000000000000000000000000001000000000000000000000000100000000000000000000,
		104'b00000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000000001,
		104'b00000000000000010001000000000001000100000000000000000000000000000000000100000000000000100000000000000000,
		104'b00000000000000000000000000000000001000000001000100000001000000000000000000000001000000000000000000000001,
		104'b00000000000000000000000000000000000000000000000000000000000100000000000100000000000100010000000000000000,
		104'b00000000000000010000000000000000000000000000000100010000000000010000000000000000000000000000000000000000,
		104'b00000000000000000000000000000001000000000000000000000001000000000000000000000001000000010000000000000001,
		104'b00000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001,
		104'b00000001000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000001,
		104'b00000000000000000000000000010000000000000000000000100010000000000000000000000001000000100000000000000010,
		104'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000010000000100000001000000000000000000000000000000000000000000000000000000000001,
		104'b00000000000000000000000100000000000000000000000100000000000100000000000000000000000000000001000100000000,
		104'b00000000000000000000000000010000000100000000000000000000000000000000000000000001000000010000000000000001,
		104'b00000000000000000000000100010000000000000000000000010000000000000000000100000000000000010001000000000000,
		104'b00000000000000000000000000010000000000000000000100000000000100000000000000010000000000010000000000000000,
		104'b00000000000000000000000000000000000100000000000000000000000100000000000000000000000000010000000000000001,
		104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000,
		104'b00000000000000000000000000010000000000000000000000000001000000000000000100000000000000010000000000000000,
		104'b00000000000000000000000000100000000100000000000100110000000100000000001000000000000000010000000000000010,
		104'b00000000000000000000000000010000000100000000000000010000000000000000000000000000000000100000000100000000,
		104'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010001,
		104'b00000000000000000000000100010001000000000000000000000001000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000010001000100000000000100000000000000000000000000000000000000010000000000000000,
		104'b00000000000000000001000000010000000100000000000000000000000100000000000000000000000000010000000000000001,
		104'b00000000000000000000000000010001000000000000000100010010000000000000000000000000000000010000000100000000,
		104'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000010001000000000001,
		104'b00000000000000000001000000010000000000000001000100010001000100000000000000000000000000110001000000000000,
		104'b00000000000000000000000000010000001000000001000100000000000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000000000000000000000000000100000000000000000000000000000000001000000000000000000000,
		104'b00000000000000000000000000000000000100000000000000000010000000000000000000000000000000100000000000010000,
		104'b00000000000000000000000000010001000000000000000000000000000100000000000100000000000000010001000000000001,
		104'b00000000000000000000000000000000000000000000000000010000000100000000000100000000000000010000000000000000,
		104'b00000000000000000000000000010001000100000000000000000001000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000000000000000100000000000100000000000000000000000000000000000100100000000000010000,
		104'b00000000000000000000000000010001000000000000000100000000000100000000000000010000000000010000000000000000,
		104'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000000000,
		104'b00000000000000000000000000000001000000000000000000010000000000000000000000000000000000010001000000000000,
		104'b00000000000000000000000000010000000100000000000000000000000000000000000100010001000000000000000000000000,
		104'b00000001000000000000000000010000000000000001000000000000000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000100000001000000000000000000000000000000000000000000000000000000100000000100010001,
		104'b00000000000000000000000000000000000000000000000100000000001000000000000000000000000000000000000100000001,
		104'b00000000000000000000000000010001000000000000000100000000000000000000000000010000000000010000000000000000,
		104'b00000000000000000000000100000001000000000000000000010000000000000000000100000001000000000000000000000000,
		104'b00000000000000000000000100010010000100000000000000000000000100000000000000000000000000010000000000000000,
		104'b00000000000000000000000000000000000000000000000100000000000000000000000100000000001000010000000100000000,
		104'b00000000000000000000000100010000000000000000000100010000000000000000000100000000000000010001000100000001,
		104'b00000000000000000000000000010000000000000000000100100000000100000000000100000000000000000000000000000010,
		104'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000001,
		104'b00000000000000000000000000000001000000000000000000010000000000000000000100000001000000010001000000000000,
		104'b00000000000000000000000000010000000000000000000000000000000000010000000000000000000000010000000000000001,
		104'b00000000000000000000000000010001000000000001000100000000000000000000000000000000000000010001000000000000,
		104'b00000000000000000000000000100000000100000000000000100000000000000000000100000000000000100000000000000000,
		104'b00000000000000000000000000000010000100000000000000000000000000000000000000000000000000010010000000000001,
		104'b00000001000000000000000100010000000000000000000100010010000000000000000100000000000000000000000100000000,
		104'b00000000000000010000000000010000000000000000000000010000000000000000001000010000000000000000000000000000,
		104'b00000000000000000000000000100010000000000000000000000000000000000000000000000000000000010000000000000001,
		104'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000010,
		104'b00000000000000010000000000010000000000000000000000010000000000000000000000000000000000000000000000000001,
		104'b00000000000000000000000000000000000000000001000100010000000000000000000000010000000000010000000000000000,
		104'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000010000000000000,
		104'b00000000000000000000000000000001000000000010000000010000000000000000001000010001000000000000000000000000,
		104'b00000000000000000001000000000001001000000000000000000000000000000000000000000000000000110001000000000000,
		104'b00000000000000000000000100010001000000000000000000000000000000000001000000000000000000010000000100010000,
		104'b00000000000000010000000000010000000000000000000000010000000000000000000000000000000000110000000000010000,
		104'b00000000000000000000000100000000000100000000000100000001000000000000000000000000000100000000000000000000,
		104'b00000001000000000000000000000000000000000000000000000001000100000000000100000000000100000000000000000001,
		104'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000100010000000100000000000000000001000000000000000000000000,
		104'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000010001000000010001,
		104'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000010001000100000000,
		104'b00000000000000010000000000000001000000000000000100000000000000000000000000010000000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000001000000000000000000000000000000010000000000000000000000000000000000100000000000000000,
		104'b00000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000100010001,
		104'b00000000000000000000000000000000000000000000000000000000000000010000000000010000000000010000001000000000,
		104'b00000000000000000000000000000001000000000001000000000000000100000000000100000000000000010000000100000001,
		104'b00000000000000000000000000000001000100000001000000000000000000000000000100000000000000010000000100000000,
		104'b00000000000000010000000000010001000000000000000000000000000000000000000100000000000000100000000000010000,
		104'b00000000000100000000000000000000000000000000000000010000000000000000000100000000000000010001000000000000,
		104'b00000000000000000000000000000000000000000000000000010000000000000000000100000001000000010000000000010000,
		104'b00000000000000010000000000000000000000000000000100010001000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000100000000000000000000000000000001000000000000000000010000000000000000000100000000,
		104'b00000000000000000000000000000001000000000000000000010000000000000000000100000001000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000000000000000100000000000100000000000100010000000000000000,
		104'b00000000000000000000000000000000000000000000000000010000000100010000000100000000000000000000000000000000,
		104'b00000000000000000000000000000000000000000001000100010000000000000000000000000000000000010000000000000000,
		104'b00000001000000000000000000010000000000000000000100000000000000000000000000000000000000000001000000000001,
		104'b00000001000000000000000000010000000000000000001000010000000100000000000000010001000000010000000100000000,
		104'b00000000000000000000000100010001000000000000000100000000000000000000000000010000000000000000000000000000,
		104'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000010000000100000001,
		104'b00000000000000000000000000010000000100000001000100000000000000000001000000000000000000010000000100000000,
		104'b00000000000000000000000000000001000000000000000000000001000000000000000000000000000000010000000000000001,
		104'b00000000000000000000000000000001000000000001000000000000000000000000000000000001000000010000000000000001,
		104'b00000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000,
		104'b00000000000000000001000000000001000100000000000100010000000000000000000100000000000000010000000000000000,
		104'b00000000000000000000000000010001000000000000000100010000000000000000000100000000000000010000000100000000,
		104'b00000000000000010000000000000000000000000000000100010000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000100000000000000000000000100010000000000000000000000000000000100000001000000000000,
		104'b00000000000000000000000000010010000100000001000100000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000100000001000000000000000100000000000000000000000000010000000000010000000000000000,
		104'b00000000000000000000000000010000000100000000000000000000000100000000000000000000000000100001000000000001,
		104'b00000001000000000000000100010001000100000000000000000000000000000000000100000000000000010000000100000000,
		104'b00000000000000000000000000010000000000000000000100000000000000000000000000010000000000000000000000010000,
		104'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000,
		104'b00000001000000000000000100010000000000000000000100010000000000000000000000000000000000000000000100000000,
		104'b00000000000000000000000000000000000100000000000000010001000000000000000100000000000000010000000100000010,
		104'b00000000000000000000000000010000000000000001001000000000000000000000000000010000000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000000000001000000000000000000000001000000010000000000000001,
		104'b00000000000000000000000000000001000100000000000000000010000000000000000000000000000000100000000000010000,
		104'b00000000000000010000000000000000000100000001000100000000000000000000000000000000000000010000000000000000,
		104'b00000000000000010000000000000000000000000000000000000000000100000000000100010000000000010000000000000000,
		104'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000100000001,
		104'b00000000000000010000000000010000000100000000000100010000000000010000000000000000000000010000000000000000,
		104'b00000000000000010000000000000000000000000000000100010000000000000000000000000000000000000001000000000000,
		104'b00000000000000000000000100010000000100000001000100000001000000000000000000000000000000010000000100000000,
		104'b00000001000000000000000000010011000000000000000000000001000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000000010000000100000000000000000000000000000000000000010000000000100000000000000000,
		104'b00000000000000000000000000100000000000000000000100000000000100000000000000000000000000000000000000000001,
		104'b00000000000000000000000000000000000000000001000000000000000100000000000000000000000000010000000100000001,
		104'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000010001000000000000,
		104'b00000000000000010000000000000000000000000000001000010000001000000000000100000001000100000000000000000000,
		104'b00000000000000010000000000000000000000000000001000010000000100000000000000000000000000000010000000000001,
		104'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000000000001000000000000000100010000000000000000000000000000,
		104'b00000000000000010000000100100000000000000000000100000000000000000000000100010000000000000000000000000000,
		104'b00000000000000000000000000000000000100000001000000000000000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000010000001000000001,
		104'b00000000000000000000000000010000000000000000000000010000000000010000000100010000000000000000000000000000,
		104'b00000000000000000000000000010000000100000000000100010000000000000000000000010000000000000000000000000000,
		104'b00000000000000000000000100000010001000000000000100000000000000000000000000000000000000100000000100000000,
		104'b00000000000000000000000100010000001000000000000000010000000000000000000000000000000000010000000100000000,
		104'b00000000000000000000000000010010000000000001000100000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000000000000000000000000000100000001000000000000000000010000,
		104'b00000000000000000000000000000000000000000000000000000001000000000000000100000000000000010001000000000001,
		104'b00000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000001,
		104'b00000000000000000000000000010000000100000000001000010000000100000000000000000000000000000000000100000000,
		104'b00000000000000010000000000010000000100000000000000000000000000000000000000000000000000010000000000000001,
		104'b00000001000000000000000000010001000100000000000100000000000000000000000100010000000000000000000000000000,
		104'b00000000000000000000000100010001000100000001000000000000000000000000000100000000000000010000000100000000,
		104'b00010000000000000000000000000001000000000000000000000000000000000000000100000000000000010000000000000000,
		104'b00000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000001,
		104'b00000000000000000000000000000001000100000001000100010000000100000000000000000000000000010000000000000001,
		104'b00000000000000000000000000000001000000000000000000010000000000000000000100000000000000010000000100000000,
		104'b00000000000000000000000100000000000000000000000000100000000100000000001000000001000000000001000100000000,
		104'b00000000000000000000000100000000000000000000000000000000000000000000000100000001000000010001000000000000,
		104'b00000000000000000000000000000001000000000001000100000000000000000000000000010000000000000000000000000000,
		104'b00000001000000000000000000010000001000000000000100000000000000000000000100000000000000010001000100000000,
		104'b00000000000000000000000000000000000100000000000100000000000000000000000000000000000000000001000000010001,
		104'b00000000000000000000000000010000000000000000001000010000000100000000000100000000000000000000000100000001,
		104'b00000000000000000000000000000000000000000000000000010000000000000000000000010001000000010000000100000001,
		104'b00000000000000010000000000010000000000000000000000000000000000000000000100010000000000010000000000000000,
		104'b00000000000100000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000000000001000000000000000000000001001000000000000000000000000000000000000000000001,
		104'b00000000000000000000000000010000000100000000000000010000000000000000000100000001000000000000000000000001,
		104'b00000000000000000000000000010000000100000000000000000000000000000000000000000000000000010000000000000001,
		104'b00000000000000000001000000010000000100000000000100100001000000000000000000000001000000100000000000000000,
		104'b00000000000000000000000000000000000100000000000000010000000100000000000100010000000000010001000100000000,
		104'b00000000000000000000000100000000000100000000000000010000000000000000000100000001000000000001000000000000,
		104'b00000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000001,
		104'b00000000000000000000000100010000001000000000000000010000000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000100100010000000000000000000010000000000000000000000000000000000010001000000000000,
		104'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000000001000000000010000100010000000000000000000100010001000000000000000000000000,
		104'b00000000000000000000000100010000000000000000000100010000000000000000000000000000000000000000001000000001,
		104'b00000000000000000000000000010001000000000000000000000001000000000000000100000000000000010000000000000000,
		104'b00000000000000000000000000010010000000000000000000000000000000000000000100000000000000010000000000000000,
		104'b00000000000000000001000000000000000000000000000000000000001000000000000000000000000000100000000000000000,
		104'b00000000000000000000000000010000000000000000000000000000000100000000001000000001000000000001000000000001,
		104'b00000000000000000000000000000000000100000001000100000000000100000000000100000000000100010000000000000000,
		104'b00000000000000000001000100000001000100000001000100000000000000000000000100000000000000010000000000000000,
		104'b00000000000000000000000000000000000100000000000100000001000000000000000000000000000100000000000000000000,
		104'b00000000000000000001000000010001000000000000000000010000000000000000000000000000000000100000000000000000,
		104'b00000000000000000001000000000000000000000000000100000000000100000000000000000000000000010000000000000000,
		104'b00000000000000000000000000000000000000000000000100000000000100000000000000000000000000000001000000000000,
		104'b00000000000000000000000000000000000000000000000100010000000000000001000000010000000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000000010001000000000000000100000000000000000000000000000001,
		104'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000001,
		104'b00000000000000000000000100000001000100000000000100000000000000000000000000010000000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000000000001000000000000000100000001000000010000000000000001,
		104'b00000000000000000000000000100000000100000001000000010001000000000000000000000000000000100001000000000001,
		104'b00000000000000000000000000100000000000000000000000000000000100000000000100000000000000010000000000000000,
		104'b00000000000000000000000000010001000100000001000100010000000000000000001000000000000000010001000100000000,
		104'b00000000000000000000000000000000000000000000000100100000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000,
		104'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000100000001000100000000000000100000000000000000000100000000000000010000000100000001,
		104'b00000000000000000000000000010000000100000000000100010000000000000000000000010000000000010000000000000001,
		104'b00000001000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000,
		104'b00000000000000000000000000000001000000000000000000000000001000000000000000010000000000000000000000000001,
		104'b00000001000000000000000000010000001000000010000100000000000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000000000010000000000000000000000000000100000000000000000000000000000000000100000001,
		104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100000000,
		104'b00000000000000000000000000010001000000000000000000000000001000000000000100000000000000000000000000000000,
		104'b00000001000000000000000000000000000000000000000100010001000000000000000000000000000000010000000000000000,
		104'b00000001000000000000000100010000000000010000000000000000000100000000000100000000000000000000000000000001,
		104'b00000001000000000001000000000000000100000000000000000000000000000000000000000000000000100000000000000000,
		104'b00000000000000000000000000010001000000000000000000010000000100000000001000000001000000000000000000000000,
		104'b00000000000000000000000000100000000000000000000100100000000000000000000000000000000000010000000100000000,
		104'b00000001000000000000000100010000000100000000000100010000000000000000000000000000000000000000000100000000,
		104'b00000000000000000001000000010000000100000001000000000000000000000000000100000000000000010000000000000001,
		104'b00000000000000000000000000100000000000000000000000000000001000000000000100000000000000010000000000000000,
		104'b00000000000000000001000000010001000000000000000000000000000000000000001000000000000000000000000000000000,
		104'b00000000000000000001000000000001000000000000000000000000000000000000000000000000000000010000000000000001,
		104'b00000000000000000000000000010001000000000000001000000000000100000000000000000000000000000000000000000000,
		104'b00000000000000010000000000000000000000000000000100000000000100000000000000000000000000000000000000000000,
		104'b00000001000000000000000000000000000100000001000000000000000100000000000000000000000000010000000000000000,
		104'b00000000000000000000000100010001000100000000000100000001000000000000000000000000000000010000000100000000,
		104'b00000000000000000000000000000000000100000000000000000001000000000000000000000000000000110001000100010000,
		104'b00000000000000000000000000000000000100000001000100000001000000000000000000000000000000010000000100000001,
		104'b00000000000000000001000000000001000000000000000100000001000000000000000100000000000000010000000000000000,
		104'b00000000000000000000000100000000000000000000000000010000000100000000000100000000000000010001000100000000,
		104'b00000000000000000000000000000000000000000000000100000000001000000000000000000001000000100000000100000000,
		104'b00000000000000000001000100000000000000000000000000000000000100000000000000000000000000010000000000000001,
		104'b00000000000000000000000000010000000100000000000000000000000100000000000100000000000000010000000100000001,
		104'b00000001000000000000000000000000000100000000000100000000000000010000000000000000000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000001,
		104'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000001000100000001,
		104'b00000000000000000000000000000001000000000000000100000000000000000001000000000000000000000000000000010000,
		104'b00000000000000000001000000000000000100000001000100000000000000000000000100000000000000010001000000000000,
		104'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000,
		104'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000100000001000000000000,
		104'b00000000000000000000000100000001000100000000000100000000000000000000000000000000000000010000000100000000,
		104'b00000000000000000000000100010000000100000000000100000000000000000000000000010000000000000000000000000001,
		104'b00000000000000000000000000010000000100000000000000010000000000000000000100000000001000100001000000000000,
		104'b00000000000000000000000000000010000100000001000000000000000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000000000000100000000000000010000000100000000000000000000000000010000000000000001,
		104'b00000000000000000000000000000001000000000000000000000000000100000000000000000000000000010000000000000001,
		104'b00000000000000000000000100000000000100000000000100010000000000000000000000000000000000000001000000000001,
		104'b00000000000000000000000000010000000100000001000000010000000000000000000100000000000000000000000000000000,
		104'b00000000000000000000000100000001000100000000000100000000000000000000000000000000000000010000000100000000,
		104'b00000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000010000,
		104'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000100000011,
		104'b00000000000000000000000000000010000100000001000100000000000000000000000000000000000000010000000100000000,
		104'b00000000000000000000000000010000000000000000000000010000000000000000000000000000000000100000000000000000,
		104'b00000000000000000000000000000000000100000000001000000001000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000010001000000000000000100000000000000010000000000000000000000000000000100000000,
		104'b00000000000000000000000000010000000100000000000000100000000000000000001000000001000000000000000000000001,
		104'b00000000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000,
		104'b00000000000000000000000000010000000100000000000000000000000000000000000100000000000000010001000100000000,
		104'b00000000000000000000000000010000000000000001000100010000000000000000000100000000000000000000000000000000,
		104'b00000000000000000000000000000000000000000000000100010000000000000001000100000000000000000000000000000000,
		104'b00000000000000000000000000000001000000000000000000010000000000000000000100000000000000100000001000000000,
		104'b00000000000000000000000000000000000000000000000000010001000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000000010001000100000000000100000000000000000000000100000001000000100000000100000001,
		104'b00000000000000000001000000000000000000000000000000010000000000000000000000000000000000010010000100000010,
		104'b00000000000000010000000000010001000000000000000000000000000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000000000010000000000000000000000000000100000000000000000000000000010000000000000001,
		104'b00000000000000000000000000000000000000000000001000000000000100010000000000000000000000000000000000000000,
		104'b00000000000000000000000000000001000000000000000000010000000100000000000100010001000000010000000000000000,
		104'b00000000000000000000000000010000000000000000000000000000000100000000000000000000000100010000000000000000,
		104'b00000000000000000000000000010000000000000000000000000001000000000000000000000000000000010000000000000001,
		104'b00000000000000000000000000100001000000000000000000000000000000000000000000000000000000100000000000000001,
		104'b00000000000100000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000,
		104'b00000000000000000000000000010001000000000000001000100000000000000000001000000000000000000001000100000000,
		104'b00000000000000000000000000010001000000000000000000000000000100000000000000000000000000100000000100000000,
		104'b00000000000000100000000000000001000000000000000100010000000000000000000100000000000000000001000000000000,
		104'b00000000000000000000000000010001000000000001001000000000000000000000000000010000000000000000000000000000,
		104'b00000001000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001,
		104'b00000000000000000000000000010000000100000000000000000000000000000000000000010000000000010001000000000001,
		104'b00000000000000010000000000000000000000000000000000000000000000010000000000000000000000100000000000000000,
		104'b00000001000000000000000000010000000100000000000100000000000000000000000000000001000000010000000100000001,
		104'b00000000000000000000000000010000000000000000000100010000000000000000000000000000000000010000000000000000,
		104'b00000000000000000001000000000000000000000000000000000000000100000000000100000000000000010000000000000000,
		104'b00000000000000000000000000000000000100000000000000000000000100000000000000000001000000010000000000000001,
		104'b00000001000000000000000000000000000100000000000000000000001000000000000000000001000000010000000000000001,
		104'b00000000000000000000000000010000000000000000000000000000000100000000000000000000000000010000000000010001,
		104'b00000000000000000000000000010001001000000000000000000000000000000000000100000001000000100000000000000000,
		104'b00000000000000010001000000000000000100000000000100000000000000000000000000010000000000100000000000000000,
		104'b00000000000000000000000100000000000000000000000000010000000000000001000000000000000000010000000000000000,
		104'b00000000000000000000000000010000000100000000001000000000000000000000000000000000000000010000000100010000,
		104'b00000000000000000001000000000000000100000000000100010001000000000000000000000000000000100000000000010000,
		104'b00000000000000000000000000010000000100000000000000000001000000010000000000000000000000010000000000000001,
		104'b00000001000000000000000000000000001000000000000000000000000100000000000100000000000000000000000000010001,
		104'b00000001000000000000000000000000000100000000000000000000001000000000000000000000000000010000000000000001,
		104'b00000000000000000000000000010000000000000000000100010000000000000000000100000000000000000000000100000001,
		104'b00000000000000000000000000100001000100000000000000000000000000000000000000000000000000000000000000000001,
		104'b00000000000000000000000000000010000100000000000000000000000000000000000100000000000000100000000000000000,
		104'b00000000000000000000000000000000000000000000000100000001000100000000000000000000000000010001000000000000,
		104'b00000000000000000000000100010001000100000000000000000000000000000000000000000000000100100000000000000001,
		104'b00000000000000000000000000000000000100000000000000000000000000000000000100000000000000000000000000000001,
		104'b00000001000000000000000100010001000100000000000000010000000000000000000100000000000000000001000000000000,
		104'b00000000000000000000000000000000000000000001000000010000000100000000000000000000000000000000000000000001,
		104'b00000000000000000000000100000000000000000000000000010001000000000000000000010000000000000000000000000001,
		104'b00000000000000000001000000000000000100000001000100000000000000000000000100000000000000010010000000000000,
		104'b00000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000,
		104'b00000001000000000000000000000001000000000000000000000000000000000000000000000000000000010000000000000000,
		104'b00000000000000000000000100000000001000010000000000000000000000000000000100000000000000100001000000000000,
		104'b00000000000000000000000000000001000000000000000100010000000000000000000000000000000000010001000100000000,
		104'b00000000000000000000000000010000000000000000000100000000000000000000000000010000000000000000000000000000,
		104'b00000000000000000000000000000011000100000000000100000000000000000000000100000000000000100000001000000001,
		104'b00000000000000000000000000010001000000000000000100000000000000000000000000000000000000000000000100000000,
		104'b00000000000000000001000000000000000000000000000100000001000000000000000100000000000000010000000000000000,
		104'b00000000000000000000000100000001000100000000000100000001000000000000000000000000000100000000000000000000,
		104'b00000000000000000000000000000000000100000000000000000001000000000000000000010000000000000000000100000001,
		104'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001,
		104'b00000000000000000000000000010001000100000001000000000001000000000000000000000000000000110000000000010000,
		104'b00000000000000000000000000100000000100000000000000000000000000000000000000000000000000100000000000010000,
		104'b00000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001,
		104'b00000000000000000000000100010010000000010000000100010000000000000000000100000000000000010000000000000000,
		104'b00000001000000000000000100000000000000000000000000000000000100000001000000000000000000000000000000000000,
		104'b00000001000000000000000000000000000000000000001000000000000000000000000000010000000000000000000000000001
	};
	
	localparam bit [7:0] alphabet [0:25] = '{
		8'b00000010,
		8'b00000011,
		8'b00000100,
		8'b00000101,
		8'b00000110,
		8'b00000111,
		8'b00001000,
		8'b00001001,
		8'b00001010,
		8'b00001011,
		8'b00001100,
		8'b00001101,
		8'b00001110,
		8'b00001111,
		8'b00010000,
		8'b00010001,
		8'b00010010,
		8'b00010011,
		8'b00010100,
		8'b00010101,
		8'b00010110,
		8'b00010111,
		8'b00011000,
		8'b00011001,
		8'b00011010,
		8'b00011011
	};
	
	// local parameters
	localparam S_IDLE      = 3'd0;
	localparam S_PRE_CALC  = 3'd1;
	localparam S_CALC      = 3'd2;
	localparam S_POST_CALC = 3'd3;
	localparam S_DONE      = 3'd4;
	
	// logics
	logic [2:0] state_r, state_w;
	logic finish_r, finish_w;
	logic [COUNT_SIZE - 1:0] word_count_r, word_count_w;
	logic [119:0] word_r, word_w;
	logic         similarity_word_w  [0:COUNT_DICT_SIZE - 1], similarity_word_r  [0:COUNT_DICT_SIZE - 1];
	logic [4:0]   similarity_value_w [0:COUNT_DICT_SIZE - 1], similarity_value_r [0:COUNT_DICT_SIZE - 1];
	logic [4:0]   max_similarity_value_r, max_similarity_value_w;
	logic [8:0]   wd_r, wd_w;
	logic [4:0]   ptr_r, ptr_w;
	
	integer i, ptr_word;
	
	// assign values
	assign o_similarity_finish = finish_r;
	assign o_similarity_word = similarity_word_r;
	
	always_comb begin
		state_w = state_r;
		finish_w = finish_r;
		word_count_w = word_count_r;
		word_w = word_r;
		similarity_word_w = similarity_word_r;
		similarity_value_w = similarity_value_r;
		max_similarity_value_w = max_similarity_value_r;
		wd_w = wd_r;
		ptr_w = ptr_r;
		
		case (state_r)
			S_IDLE: begin
				finish_w = 1'b0;
				if (i_similarity_start) begin
					state_w = S_PRE_CALC;
				end
			end
			S_PRE_CALC: begin
				// calculate word count
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[0] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[1] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[2] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[3] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[4] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[5] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[6] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[7] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[8] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[9] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[10] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[11] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[12] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[13] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[14] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[15] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[16] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[17] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[18] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[19] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[20] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[21] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[22] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[23] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[24] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
					end
				end
				for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 8) begin
					if (alphabet[25] == i_similarity_word[ptr_word +: 7]) begin
						word_count_w = word_count_w + 104'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
					end
				end
				
				state_w = S_CALC;
			end
			S_CALC: begin
				// calculate each similarity value
				if (wd_r == COUNT_DICT_SIZE - 1) begin
					state_w = S_POST_CALC;
				end else begin
					for (ptr_word = 0; ptr_word < 120; ptr_word = ptr_word + 4) begin
						// output the smaller value
						if (count_dict[wd_r][ptr_word +:3] >= word_count_r[ptr_word +:3]) begin
							similarity_value_w[wd_r] = similarity_value_w[wd_r] + {100'b0, word_count_r[ptr_word +:3]};
						end else begin
							similarity_value_w[wd_r] = similarity_value_w[wd_r] + {100'b0, count_dict[wd_r][ptr_word +:3]};
						end
					end
					
					if (similarity_value_w[wd_r] >= max_similarity_value_r) begin
						max_similarity_value_w = similarity_value_w[wd_r];
					end
					wd_w = wd_r + 1;
				end
			end
			S_POST_CALC: begin
				// find the biggest 20 values
				if (ptr_r >= 20) begin
					state_w = S_DONE;
				end else begin
					for (ptr_word = 0; ptr_word < COUNT_DICT_SIZE; ptr_word = ptr_word + 1) begin
						if (ptr_w >= 20) begin
							break;
						end
						if (similarity_value_w[ptr_word] == max_similarity_value_r) begin
							similarity_word_w[ptr_word] = 1'b1;
							ptr_w = ptr_w + 1;
						end
					end
				end
				
				max_similarity_value_w = max_similarity_value_r - 5'd1;
			end
			S_DONE: begin
				finish_w = 1'b1;
				state_w = S_IDLE;
			end
		endcase
		
	end

	always_ff @ (posedge i_similarity_clk or posedge i_similarity_rst_n) begin
		if (i_similarity_rst_n) begin
			state_r                <= S_IDLE;
			finish_r               <= 1'b0;
			word_count_r           <= 104'b0;
			word_r                 <= 120'b0;
			similarity_word_r      <= '{500{1'b0}};
			similarity_value_r     <= '{500{5'b0}};
			max_similarity_value_r <= 5'b0;
			wd_r                   <= 9'b0;
			ptr_r                  <= 5'b0;
		end else begin
			state_r                <= state_w;
			finish_r               <= finish_w;
			word_count_r           <= word_count_w;
			word_r                 <= word_w;
			similarity_word_r      <= similarity_word_w;
			similarity_value_r     <= similarity_value_w;
			max_similarity_value_r <= max_similarity_value_w;
			wd_r                   <= wd_w;
			ptr_r                  <= ptr_w;
		end
	end
endmodule

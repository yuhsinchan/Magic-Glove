module Similarity(
	input          i_similarity_clk,
	input          i_similarity_rst_n,
	input          i_similarity_start,
	input [119:0]  i_similarity_word,
	output         o_similarity_finish,
	output[9:0]    o_similarity_word[0:19]
);

	parameter COUNT_DICT_SIZE = 600;
	parameter COUNT_SIZE = 26 * 4;

	localparam bit [COUNT_SIZE - 1:0] count_dict [0:COUNT_DICT_SIZE - 1] = '{
        104'b00000000000100000000000000010000000000000000000000010000000000000000000000000000000000010000000000000000,
        104'b00000001000000000000000000010000000100000000000000010000000100000000000000000000000000100000000100000000,
        104'b00000000000000000000000100000000000100000010000000000000000100000000000000000000000000010000000000000000,
        104'b00000000000000000000000100010000000100000000000100010000000000000000000000000000000100100000000000000000,
        104'b00000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000,
        104'b00000001000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000,
        104'b00000000000000000000000100000000000000000000000000000000000100000000000000000000000100000000000000000000,
        104'b00000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000,
        104'b00000000000000000000000100000000000100000000000000000000000000000000000000000000000000010001000000000000,
        104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000000000001,
        104'b00000000000000000000000100000000000000000000000000000000000100010000000000000000000000000000000100000000,
        104'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000,
        104'b00000000000000000001000000000000000100000000000000000000000000000000000000000000000100100000000000000000,
        104'b00000000000000010000000000000000000100000000000100010000000000000000000000000000000000000000000000010000,
        104'b00000000000000000000000000010000000000000000000000010000000000010000000000010000000000000000000000000001,
        104'b00000000000000000000000100000010000000000010000100000000000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000100000001,
        104'b00000001000000000000000000100000000100000001000000000000000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000000000000000000000010000100000000000100000000000000000000000000100000000000000000,
        104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000000010000,
        104'b00000000000000000000000000000000000000000000000100000000000100000000000000010000000000000001000000000000,
        104'b00000000000000000000000000010001000000000000000100000000000000000000000000000000000000000000000100000000,
        104'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000001,
        104'b00000000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000000,
        104'b00000000000000000000000000000001000100000001000000000000000000000000000000000001000000010001000000000001,
        104'b00000000000000000000000000000001000000000000000000000000000100000000000000000000000000100000000000000000,
        104'b00000000000000000000000000010000001000000000000100000000000000000000000000010000000000010000000000010000,
        104'b00000000000000000000001000000011000000000000000000000000000100000000000000000000000100010000001000000000,
        104'b00000000000000000000000000000000000000000000001000000000000100000000000000000000000100000000000000000000,
        104'b00000000000000000000000100000001000000000000000000010000000000000000000000010000000000000001000000010001,
        104'b00000000000000000000000000000001000000000000000000000001000000010000000000000000000000010000000000000001,
        104'b00000000000000000000000000000000000100000000000100000000000000000000000000000000000000000000000000000000,
        104'b00000000000000000000000000000000000100000000000000000000000000000000000000010000000000100000000100000000,
        104'b00000000000000000000000000000000000000000000000000000000000100000000000000000001000000010000000000000000,
        104'b00000000000000000000000000010001000000000000000100000000000100000000000000010000000000010000000100000000,
        104'b00000000000000000000000100000001000000000000000000000000000000000000000000010000000000000000000100000000,
        104'b00000001000000000000000100000000000000000000000000000000000100010000000000000000000000000000000100000000,
        104'b00000000000000000000000000000000000000000000000000000000000100000000000000000001000000000001000000000001,
        104'b00000000000000010000000000000000000000000000000100000001000100000000000000000000000000100000000100000000,
        104'b00000000000000000000000000000000000000000000000000010000000000000000000000010000000000000001000000000001,
        104'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000010000000000000001,
        104'b00000000000000000000000000000001000000000000000100000001000000000000000000000000000000010000000100000000,
        104'b00000000000000000000000000010001000100000000000100000000000000000000000000010000000000010000000000000000,
        104'b00000000000000000000000000000000000000000000000100010000000000000000000000000000000000010000000100000000,
        104'b00000001000000000000000000010001000100000000000100000000000000000000000000000000000000000000000000000000,
        104'b00000000000000000001000000000000000100000000000000000000000100000000000000000000000000100000000100000000,
        104'b00000000000000000000000000000000000100000001000100000000000000010000000000000000000000000000000000000000,
        104'b00000000000000000000000000000010000100000000000100000000000000000000000000000000000000000000000100000001,
        104'b00000000000000000001000000000000000100000000000000010000000000000000000000000000000000100000000000000000,
        104'b00000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000001,
        104'b00000000000000000000000000010000000100000000000100000001000000000000000000010000000000010000000000000000,
        104'b00000000000000000000000000000000000100000000000100000000000000000000000000000000000000000001000000000001,
        104'b00000000000000000000000000000001000000000000001000010001000000000000000000000000000000100000000000000000,
        104'b00000001000000000000000000100000000000000000000100000000001000000000000000000000000000000000000000000001,
        104'b00000001000000010000000000100000000000000000000000010000000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000100000000000000000000000000000001000100000000000000010000000000010000000000010000,
        104'b00000000000000000000001000000001000100000000001000000001000000000000000000010000000000000000000000000000,
        104'b00000000000000010000000000000000000100000000000100000000000100000000000000000000000000000001000000000000,
        104'b00000000000000000000000000000001000000000001000100000000000000010000000000000000000000010000000000000000,
        104'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000100100000000000000000,
        104'b00000000000000010000000000000000000000000000000000000000001000000000000000000000000000000000000000000001,
        104'b00000000000000000000000000000000000000000000000000010000000000000000000000010000000000010000001000000001,
        104'b00000000000000000000000100010001000000000000000100010000000000000000000000010000000000000001000000000001,
        104'b00000000000000000000000000000000000100000000000100100000000000000000000000000000000000100001001000000000,
        104'b00000000000000000000000000000000000100000000000000000000000000000000000000000001000000010000000100000001,
        104'b00000000000000000000000000000010000100000000000000000000000100000000000000000000000000100000000100000001,
        104'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000,
        104'b00000000000000000000000000010000000100000000000000010000000000000000000000000001000000110000000000000001,
        104'b00000000000000000000000000000000000000000001000000000000000000010000000000000000000000100000000000000000,
        104'b00000000000000000000000000010000000100000000000100010000000000000000000000010000000000010000000000000001,
        104'b00000000000000000000000100000000001000000000000000000001000000000000000000010001000000010000000000010001,
        104'b00000001000000010000000000010001001100000000000000000000000000000000000000000000000000010000000000010001,
        104'b00000000000000000000000000010001000000000000000000000000000100010000000000000000000000000000000000000001,
        104'b00000000000000000000000000000000000000000000000000010000000100010000000000000000000000010000000000000001,
        104'b00000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000100000001,
        104'b00000000000000010000000000000000000100000000000100000000000000000000000000000000000000000001000000000000,
        104'b00000000000000010000000000000001000000000000000100010000000000010000000000000000000000000000000000000000,
        104'b00000000000000000000000000010000000000000000000000000000000100000000000000000000000100010000000000000000,
        104'b00000000000000000000000000010000000000000001000100000001000100000000000000000000000000100001000100000000,
        104'b00000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000001,
        104'b00000000000000000000000100000001000100000000000100000000000100000000000000010000000000010001000000000000,
        104'b00000000000000000000000000010010000100000000000000000000000000000000000000000000000000100001000000000000,
        104'b00000000000000000000000000000001000000000000000000010000000000010000000000000000000000000000000100000001,
        104'b00000001000000000000000000000000000000000000000100010000000000000001000000000000000000100001000000000000,
        104'b00000000000000000000000100100000000100000000000000000000000000000000000000010000000000000000000000000000,
        104'b00000000000100000000000100000001000000000000000000000000000000000000000000000000000000100000000100000000,
        104'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000100000001,
        104'b00000000000000000000000000000000000100000001000000000000000000010000000000000000000000000000000000000001,
        104'b00000000000000000000000000010010000100000000000100000000001000000000000000000000000000000000000000000000,
        104'b00000000000000000000000100000000000000000001000000000000000000000000000000000000000000000000000100000000,
        104'b00000000000000000000000000000000001000000001000000000000000000000000000000000000000100100000000000000000,
        104'b00000000000000010000000000000000000000000000000100000000000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000000010001000000000001000100000000000000000000000000000000000000000000000000000000,
        104'b00000000000000000000000100000010000000000000000000000000000000000000000000000001000000010000000000000000,
        104'b00000000000000000000000000000010000000000000000000000000000100000000000000000000000000010000000000010000,
        104'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000000001,
        104'b00000000000000000000000100000000000000000000000100000000000100000000000000000000000000000001000100000000,
        104'b00000000000000000000000000000000000000000000000000000000000000010000000000010000000000010000001000000000,
        104'b00000001000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000000,
        104'b00000000000000000000000000000011000000000000000000000001000000000000000000000001000000100000000000000001,
        104'b00000000000000000000000000010000000000000000000100000000000000000000000000000001000000000000000000000000,
        104'b00000000000000000000000100010000000000000000000000000000000100000000000000000000000000000001000000000001,
        104'b00000000000000000000000000000001000000000000000000010000000000000000000000010000000000000001000000000001,
        104'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001,
        104'b00000000000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000001,
        104'b00000000000000000001000000000000000000000000000100000000000100000000000000000000000000010000000000000000,
        104'b00000000000000000000000000000001000000000000000000000000000100000000000000000000000000000001000000000010,
        104'b00000000000000000000000000010000000000000000000000000001000000000000000000010000000000010000000000000000,
        104'b00000000000000000000000000000000000000000000001000010000000100000000000000000000000000010001000000000000,
        104'b00000000000000000000000000000000000000000000000100010000000000000001000000010000000000000000000000000000,
        104'b00000001000000000000000000000000000000000000000100010001000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000100000000000000000000000000010000000100000000000000010000000000000000000100000000,
        104'b00000000000000000000000000000001000000000000000000010000000000000000000000000000000000100001000000000000,
        104'b00000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000000010000,
        104'b00000000000000000000001000010000000000000000000100010000000000000000000000010001000000000001000000000000,
        104'b00000000000000000000000100000000000000000000000000000000000100000000000000000000000000010000000000010000,
        104'b00000000000000000000000000100000000100000000000100000000000000000000000000010000000000000000000000000001,
        104'b00000000000000000000000000000000000000000001000000000000000100000000000000000000000000010000000100010010,
        104'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000,
        104'b00000000000000000000000000000001000000000000000000010000000000000000000000010000000000010000001000000001,
        104'b00000000000000000000000000010001000000000000000000000000000000010000000000000000000000000000000000000001,
        104'b00000000000000000000000100000000001000000000000000000000000000000000000000000001000000010000000000010000,
        104'b00000000000000000000000000000001000000000000000000010000000000000000000000000000000000100000000000000000,
        104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000,
        104'b00000000000000000000000000000000000100000000000000000000000000000000000000010000000000010001000000000001,
        104'b00000000000000000000000000100001000000000000000100010000000000000000000000000000000000010000000100000000,
        104'b00000000000000010000000000000000000000000000000000000000000000010000000000000000000000010000000000000001,
        104'b00000000000000000000000000000000000000000000000000010000000000000001000000000000000000010000000000000001,
        104'b00000000000000000000000000000000000100000000000100010000000000000000000000000001000000010000000000000001,
        104'b00000000000000000000000100100001000000000000000000010000000000000000000000000000000000010001000000000000,
        104'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000100100000000000000000,
        104'b00000000000000000000000000010000000000000000001000000000001000000000000000000000000100000000000000010001,
        104'b00000000000000010000000000000001000100000000000100000000000000000000000000000000000000000001000000000000,
        104'b00000000000000000000000000000000000000000000000100000000000000010001000000000000000000010000000000000000,
        104'b00000000000000000000000000000001000000000000000100000000000100000000000000000000000000010000000000000000,
        104'b00000000000000000000000000000000000100000000000000000000000000000000000000010000000000100000000000000000,
        104'b00000000000000000000000000000000000100000000000100000000000000000000000000000000000100000000000000000000,
        104'b00000000000000000000000000000000000100000000000000000000000000000000000000010000000000010000000000000001,
        104'b00000000000000010000000000000000000000000000000000000000000100010000000000000000000000000000000000000001,
        104'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000100000000000000000001,
        104'b00000000000000000000000100010001000000000000000000000000000000000000000000010000000000000000000000000000,
        104'b00000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000000,
        104'b00000000000000000000000000000001000100000000000000010000000100000000000000000000000000100001000000000000,
        104'b00000000000000000000000100000000000100000000000000010000000000000000000000010000000000000000000100010000,
        104'b00000000000000010000000000010001000000000000000000000000000000000000000000000000000000010000000000000001,
        104'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000100000000000000000001,
        104'b00000000000000000000000100000000000000000000000100000000000000000000000000010001000000000000000100000000,
        104'b00000001000000000000000100010001000100000000000000000000000000000000000000000000000000000001000000000010,
        104'b00000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001,
        104'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000001,
        104'b00000000000000000000000100010000000000000000000100000000000000000000000000000000000000000000000000010001,
        104'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000100000000000000000001,
        104'b00000000000000000000000000000001000000000001000000000000000100000000000000000000000000100000000000000001,
        104'b00000000000000010000000000000000000000000000000100000000000100000000000000010000000000010000000000000000,
        104'b00000000000000000000000000010000000000000000000000000000000100000000000000000000000000010000000000010000,
        104'b00000000000000000000000100000001000100000010000000000000000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000000010000000000000000000000000001000000000000000000000000000000100000000000000000,
        104'b00000001000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000001,
        104'b00000000000000000000000000010010000000000001000000000000000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000000000001000000000000000100010000000000000000000000000000000000000000000000000000,
        104'b00000000000000000000000000010000000100000000000100000000000000000000000000000001000100010000000000000000,
        104'b00000000000000010000000100000000000100000000000100010000000100000000000000000000000100010001000000000000,
        104'b00000000000000000000000100000000000000000000000000010000000000000000000000000000000100000000000000000000,
        104'b00000000000000000000000000000000000100000000000100010000000000000000000000000000000000000000000000010000,
        104'b00000000000000000000000000010000000000000000000100010000000000000000000000000000000000000000000000000000,
        104'b00000000000000000000000000000000000100000000000000010000000000000000000000000000000000010000001000000001,
        104'b00000001000000000000000000000000000000000000000100010000001000000000000000000000000000010000000000000000,
        104'b00000000000000010000000100000000000000000000000100010000000000000000000000000000000000000001000000000000,
        104'b00000000000000000000000000000000000000000000001000000000000000000000000000000001000000000001000000000000,
        104'b00000001000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000001,
        104'b00000001000000000000000000000000000000000000000100010000000100000000000000000000000000000000000000000000,
        104'b00000000000000010000000000010000000000000000000100010000000000000000000000000000000000000000000000000000,
        104'b00000000000000000000000000000000000000000000000100010001000000000000000000000001000000000000000000000001,
        104'b00000001000000000000000100000000000000000010000000010000000000000000000000010000000000000000000000000001,
        104'b00000000000000000000000000000001000000000000000000000000000000000000000000000001000000010000000000000001,
        104'b00000000000000000000000000010000000100000000001000010000000100000000000000000000000000000000000100000000,
        104'b00000000000000000000000000010001000000000000000000000000000000000000000000000000000000010000000000000001,
        104'b00000000000000000000000000000000000100000000000100000000000000000000000000000000001000000001000000000001,
        104'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000010001000000000000,
        104'b00000000000000000000000000000000000000000000000100000000000100000000000000000001000000000001000000000000,
        104'b00000000000000000000000100000000000100000000000000000000000100000000000000000000000000010000000100000000,
        104'b00000000000000000000000000010000000000000000000000000000000100000000000000100000000000010000000000000001,
        104'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000001000000000001,
        104'b00000001000000000000000100000000000100000000000100000000000000000000000000000000000000000000000000000000,
        104'b00000001000000000000000000000001000000000000000000010000000000010000000000000000000000010000000000000001,
        104'b00000001000000000000000000000000000000000000000000000000000100000000000000000000000000010010000000000001,
        104'b00000000000000000000000000000000000100000001000000000000000000000000000000000001000000010000000000000001,
        104'b00000000000000000000000000000000000000000000000000010000000100000000000000000001000000010000000000000001,
        104'b00000000000000000000000100010000000000000000000000000000000000000000000000010001000000000000000100000001,
        104'b00000001000000000000000100000000000000000000000000000000000000000000000000010000000000000000000100100000,
        104'b00000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000,
        104'b00000000000000000000000000000000000100000000000100000001000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000000010000000000000000000000010000000000000000000000000000000000010000000000000001,
        104'b00000000000000000000000000000000000100000000000100000000000000000000000000000000000100100000000000010000,
        104'b00000000000000000000000000010000001000000000000000010000000000000000000000010001000100010001000000000010,
        104'b00000001000000000000000000000001000000000000000000000000000000000000000000000000000000010000000000000001,
        104'b00000000000000000000000000010001000100000000000000000000000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000000000001000000000000001000010000000000000000000000000000000000000000000000000000,
        104'b00000000000000010000000000000000000000000000000100010000000000000000000000000000000000000000000000000000,
        104'b00000000000000000000000100000000000100000001000100000000000000000000000000000000000000000001000000000000,
        104'b00000000000000000001000000000000001000000000000100000000000000000000000000000000000000100000000100000000,
        104'b00000000000000000000000000000000000100000000000000000000000100000000000000000000000000100001000000000000,
        104'b00000001000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000,
        104'b00000000000000000000000000010001000000000000000000000000000000000000000000000000000000010000000000010000,
        104'b00000000000000000000000100000000000100000000000000000000000100000000000000000000000100010000000100000001,
        104'b00000000000000010000000000000000000000000000000100000000000000000000000000010000000000000000000000000000,
        104'b00000000000000000000000100010001001000000000000000010000000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000100000001000000000001000000000001000000000000000000000000000000000000000100000001,
        104'b00000000000000000000000000100001000000000000001000000001000000000000000000000000000000000000000000010000,
        104'b00000001000000000001000000000000000100000000000000000000000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000100010001000000000000000000000000000000000001000000000000000000000000000000000000,
        104'b00000000000000010000000000000000000000000000000100000000000000000000000000010000000000000000000000000000,
        104'b00000001000000000000000000000000000100000001000000000000000100000000000000000000000000010000000000000000,
        104'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000001,
        104'b00000000000000000000000000000000000100000000000000000000000000000000000000010001000000010001000100000001,
        104'b00000000000000000000000100000001000000000000000000000000000000000000000000000000000000010001000000000000,
        104'b00000000000000000000000000010000000100000000000000010000000000000000000000000000000000100000000000000000,
        104'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000010000000000000000,
        104'b00000000000000010000000000000001000000000000000100000000000000000000000000010000000000000000000000000000,
        104'b00000000000000000000000000000000000100000000000000010000000000000000000000000001000000100000000000000000,
        104'b00000000000000000000000000000000000000000000000100000000001000000000000000000000000000000001000000000000,
        104'b00000000000000000000000000010000000000000000000100000000000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000100110010000000000001,
        104'b00000000000000000000000000010001001000000000000000010000000000000000000000000001000000010000000000000001,
        104'b00000000000000000000000100000000000100000000000100000000000000000000000000000000000100000000000000000000,
        104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100010000000100000001,
        104'b00000000000000000000000000000001000000000001000000000000000000010000000000000000000000010000000000000001,
        104'b00000000000100000000000000010000000000000001000000000000000000000000000000000000000000100000000100000000,
        104'b00000000000000000000000000000001000100000000000100000000000000000000000000010000000000010000000000000000,
        104'b00000000000000000000000100010000000000000000000100000000000000000000000000010000000000000000000100000000,
        104'b00000000000000000000000000000001000100000000000100100000000000000000000000000001000000000001000000000001,
        104'b00000000000000000000000000010000000100000000000000000000001000000000000000000000000000010000000000000001,
        104'b00000000000000000001000000000000000000000000000000010000000100000000000000000000000000110000000000000000,
        104'b00000000000000000000000000100001000000000000000000000000000100000000000000000000000000010000000000000001,
        104'b00000000000000010000000000010000000100000000000000000000000000000000000000010000000000100000000000000001,
        104'b00000000000000000000000000010000000000000000000100000000000000000000000000010000000000000000000000010000,
        104'b00000000000000000000000000010000000000000000001000000000000100000000000000010000000000010000001000000001,
        104'b00000000000000010000000000000000000100000001000100000000000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000100010001000100000000000100000001000000000000000000000000000000010000000100000000,
        104'b00000000000000010000000000010001000100000000000100010001000100000000000000000000000000100000000000000001,
        104'b00000000000000010000000000000001000000000000000100000000000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000100000000000100000000000000000000000000000000000000000000000000010000000100000000,
        104'b00000001000000000000000000010001000000000000000000000000000000000000000000000000000000000000000000000001,
        104'b00000000000000000000000000000001000000000000000000000000000100010000000000000000000000000000000100000001,
        104'b00000000000000000000000000000001000000000000000000000001001000000000000000000000000000100001000000000000,
        104'b00000000000000010000000100000000000000000000000000000000000100000000000000000000000100000000000000000001,
        104'b00000000000000000000000000010001000100000000000000000001000000000000000000000000000000000000000000000001,
        104'b00000000000000000000000100000000000000000000000000000000001000000000000000000000000100000000000000000000,
        104'b00000000000000000001000000000000000000000000000000000000000100000000000000000000000000100000000000000001,
        104'b00000001000000000000000000000000000000000000000000000000000100000000000000000000000000000001000000000001,
        104'b00000000000000010000000000000000000000000000000100010000000000000000000000000000000000000001000000000000,
        104'b00000000000000000000000000010001000100000000000100000000000000000000000000000000000000000000000000000000,
        104'b00000000000000000000000100000001000100000000000000000000000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000000000000000000000000000000010001000000000000000000000000000000010000000000000001,
        104'b00000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000010000,
        104'b00000000000000000000000100010000000100000000000000000000000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000100010000000000000000000100010000000000000000000000000000000000000000000100000000,
        104'b00000000000000000000000000000000000100000000000000010000000000000000000000000001000000010001000000000001,
        104'b00000000000000010000000000000000000100000000000000000000000000000000000000010000000000100000000000000000,
        104'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001,
        104'b00000000000000000000000000010001000000000000000100000001000000000000000000000000000000010001000000000000,
        104'b00000000000000000000000100010000000000000000000100000001000000000000000000010000000000000000000000000000,
        104'b00000000000000000000000000010000001000000000000000000000000000000000000000000001000000100000000000000000,
        104'b00000000000000000000000000000010000000000001000000000000000000000000000000000000000000000000000000000001,
        104'b00000001000000000000000000000000000100000000000000000000000000000000000000000001000000000000000000000001,
        104'b00000000000000000000000000000000000100000000001000000000000100000000000000000000000000010000000100000000,
        104'b00000000000000000000000000010000000000000000000000100001000100000000000000000001000000100000000000000001,
        104'b00000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000001,
        104'b00000000000000000000000000000001000100000000000000000000000100000000000000010000000100100000000000000000,
        104'b00000000000000000000000000000000000000000000000000000000000100010000000000000000000000000000000100010001,
        104'b00000000000000000000000100000000000000000001000000000000000000000000000000000000000000000000000000000000,
        104'b00000000000000000000000100010010000000000000000000000000000000000000000000000010000000100001000000000000,
        104'b00000000000000000001000000000000000000000000000100000001000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000001,
        104'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000100000001,
        104'b00000000000000010000000000010000000100000000000100010001000100000000000000000000000000100000000000000001,
        104'b00000000000000000000000100100001001000000000000000010000000000000000000000000000000000010000000000000010,
        104'b00000000000000000000000100000000000000000000000000010000000000000000000000000001000000000000000000000000,
        104'b00000000000000000000000000010001000100000000000100000000000000000000000000010000000000000000000000000000,
        104'b00000000000000000000000000010000000100000000000000000000000000000000000000000001000000010000000000000001,
        104'b00000000000000000000000100010000000100000000000000000000000000000000000000010000000000000000000000000000,
        104'b00000000000000000000000000010001000100000000000000000000000000000000000000000000000100010000000000000001,
        104'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000001,
        104'b00000000000000000000000000010000000000000000000000000000000000000000000000000001000000010000000000000000,
        104'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000100000000000010000,
        104'b00000000000000000000000000010000000100000000000000000000000000000000000000000000000100010000000000000001,
        104'b00000000000000000000000100000010000000000000000100010000000000000000000000000000000000000001000000000000,
        104'b00000001000000010000000000000001000000000000000000000000000100000000000000000000000000000000000000000010,
        104'b00000000000000000000000100000001000000000000000000000000000000000000000000000000000000100000000100010001,
        104'b00000000000000000000000000000001000000000000000000000000000000000000000000010000000000010000000000000000,
        104'b00000000000000000000000100010000000000000000000100000000000000000000000000000000000000000001000000010000,
        104'b00000000000000000000000000010001000000000000000100000001000000000000000000100000000000010000001000000010,
        104'b00000000000000000000000000000001000100000000000000000000000000000000000000000000000000010000000000000001,
        104'b00000000000000010000000000000001000100000000000000010000000000000000000000000000000000010000000000000001,
        104'b00000000000000000000000000010001000000000000000100010000000000000000000000010000000000010000000000000000,
        104'b00000000000000000000000000000001000000000000000100010000000000000000000000000000000000010001000100000000,
        104'b00000000000000000000000100000001000000000000000000010000000000000000000000000000000000000000000000000000,
        104'b00000001000000000000000000000000000000000000000000010000000000000000000000000000000000000001000100000001,
        104'b00000000000000010000000000010000000000000000000000010000000000000000000000000000000000000000000000000001,
        104'b00000001000000000000000000000000000000000000000100000000000000000000000000000000000000000001000000010000,
        104'b00000000000000000000000100010000000000000000000000000000000000000000000000000000000000000000000100000000,
        104'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000001000000000001,
        104'b00000000000000000001000000000000000000000001000100000000000100000000000000000000000000100001000000000000,
        104'b00000000000000000000000000000000000000000001000000000000000100000000000000000000000000010000000000000001,
        104'b00000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000000001,
        104'b00000000000000000000000000000000000000000000000100010000000000000000000000000000000000010000000000010000,
        104'b00000001000000000001000000000000000000000000000100000000001000000000000000000000000000010000000000000000,
        104'b00000000000000000000000000010001000100000000000000000000000000010000000000000000000100010000000000010010,
        104'b00000000000000000000000000000001000000000000000100010000000000100000000000000000000000000000000100000000,
        104'b00000001000000000000000000010000000000000001000000010000000100000000000000000000000000010000000000000000,
        104'b00000000000000000000000000000000000000000001000000010000000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000000000010000000000000000000010000000000000000000000000000000000100000000000000000,
        104'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001,
        104'b00000001000000000000000000010000000000000000000000000000000100000000000000100000000000010000000000000001,
        104'b00000000000000000001000000000000000100000000000100000000000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010011,
        104'b00000000000000000000000000000000000000000000000100010001000000000000000000000001000000000000000000000001,
        104'b00000000000000000000000000000000000100000000000000000001000000000000000000000000000000000000000000000001,
        104'b00000000000000000000000000010000000100000000000000000000000000000000000000010000000000100000000000000000,
        104'b00000000000000000000000000000000000000000000000000000001000000000000000000000001000000010000000000000001,
        104'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000100000001,
        104'b00000001000000000001000000010001000000000000000000010000000000000000000000000000000000100000000000000000,
        104'b00000000000000010000000000000000000000000000000100010000000000000000000000000000000000010001000000000000,
        104'b00000001000000000000000000000000000000000010000000000000000000000000000000010000000000000000000000000001,
        104'b00000001000000000000000000000000000100000000000000000000000100000000000000010000000000000001000000000001,
        104'b00000000000000000000000000000010000000000000000100000000000000000000000000010000000000010000000000000000,
        104'b00000000000000000000000000010001000000000000000100000000000100000000000000000000000000000000000000000000,
        104'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000100001000100000010,
        104'b00000000000000000000000000000001000000000000000000000000000000010000000000000000000000010001000000000001,
        104'b00000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000000001,
        104'b00000001000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000,
        104'b00000000000000010000000000000000000100000000000100010000000000000000000000000000000000010001000100000000,
        104'b00000000000000000000000100000000000100000000000100000000000000000000000000010000000000000000000000000000,
        104'b00000000000000000000000000000000000000000000000000010001000000000000000000000000000000010000000000000000,
        104'b00000000000000010000000000010000000000000000000000010000000000000000000000000000000000110000000000010000,
        104'b00000000000000010000000000010000000000000000000000010000000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000100000001000000000001000100000000000000000000000000000000000000000000000000000000,
        104'b00000000000000000000000000010000001000000000000000000000000000000000000000010000000000010000000000000001,
        104'b00000000000000000000000000000000000000000000000100000000000000000000000000000001000000000001000000000000,
        104'b00000000000000000000000000010001000000000000000100000000000000000000000000010000000000000000000000000000,
        104'b00000001000000010000000000000000000000000000000100000000001000000000000000000000000000010000000000000000,
        104'b00000001000000000000000100010000000000000000000000010000000000000000000000010001000000000000000000000001,
        104'b00000001000000000000000100010000000000000000000100000000000000000000000000010000000000000000000000000000,
        104'b00000000000000000000000000000000000100000000000100000001000000000000000000000000000100000000000000000000,
        104'b00000000000000000000000000010001000100000000000100010000000000000000000000000001000000000000000000000000,
        104'b00000001000000010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000,
        104'b00000001000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000,
        104'b00000000000000000000000000000000000000000000000100000000000100000000000000000000000000000001000000000000,
        104'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000001,
        104'b00000000000000000000000000000000001000000000000000000001000100010000000000000000000000100000000000010010,
        104'b00000000000000010000000000000000000000000000000100010000000000000000000000000000000000000000000000000000,
        104'b00000000000000000000000000000010000000000000000100000001000000010000000000000000000000010000000000000000,
        104'b00000000000000010000000000000000000000000000000100010000000000000000000000000000000000000000000000000000,
        104'b00000001000000010000000000000000000100000000000000000000000100000000000000000000000000010000000000000001,
        104'b00000010000000000000000000010001000100000000000000000000000000000000000000000000000000100001000000000001,
        104'b00000000000000000000000100000001000000000001000000000000000000000000000000000000000000010001000000000001,
        104'b00000000000000000000000000010000000000000000000100000000000100000000000000000000000000000001000000000000,
        104'b00000001000000000000000000000001000000000000000000000000000000000000000000000000000000100000000000000000,
        104'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000010000000100000001,
        104'b00000001000000000000000000000001000000000000000000000000000100000000000000000000000000000001000000000001,
        104'b00000000000000000000000000010000000100000000000000000000000000000000000000010000000000010000000000000001,
        104'b00000000000000010000000000000000000000000000000000000000001000000000000000000000000000010000000000000000,
        104'b00000000000000000000000000010000000100000001000000010000000000000000000000000000000000010000000000000001,
        104'b00000000000000000000000000100000000100000000000000000000000000000000000000000000000000010000000000000001,
        104'b00000000000000000000000000010000000000000000000000000000000000000000000000010000000000010000000000000000,
        104'b00000000000000010000000000000001000000000000000100000000000100000000000000000000000000000000000000000000,
        104'b00000000000000000000000000000000000000000000001000000000000100000000000000000000000000000000000100000000,
        104'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000010001000000010001,
        104'b00000000000000010000000000000000000100000000000100000000000000010000000000000000000000000000000000000000,
        104'b00000000000000000000000000010001000000000000000000000000000000010000000000000000000000010000000000000001,
        104'b00000000000000000000000000000001000000000001000000000000000100000000000000000000000000100000000000000000,
        104'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000010001000000000001,
        104'b00000000000000000001000100000001000100000000000100010000000000000000000000000000000000010000000000000000,
        104'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001,
        104'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000010001000000000001,
        104'b00000000000000000000000000010001000000000000000100000000000000000000000000010000000000010000000000000000,
        104'b00000000000000000000000000000000000000000000000000000001000100000000000000000000000000010000000000000001,
        104'b00000000000000000000000000010001000100000000000000000001000000000000000000000000000000010000000000000001,
        104'b00000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000001,
        104'b00000001000000000000000000000000000100000000000100000000000000010000000000000000000000000000000000000000,
        104'b00000000000000000000000000000000000000000000000100000000000000000000000000000001000000000001000000000000,
        104'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000010001000000000000,
        104'b00000000000000000000000000000000000000000000000100010000000100000000000000000000000000010000000000000001,
        104'b00000001000000000000000000000001000000000000000000000000001000000000000000000000000000000000000000000001,
        104'b00000000000000000000000000000000000000000000000100000001000000000000000000000000000000010000000100000000,
        104'b00000000000000000000000000000000000100000000000000000000000100000000000000000001000000010000000000000001,
        104'b00000000000000000000000100000000000100000000000000010000000000000000000000000000000000010001000000000000,
        104'b00000000000000000000000000010001000000000000000000000000000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000000100000000100000000000000000000000000000000000000000000000000100000000000010000,
        104'b00000000000000000000000100000001000000000000000100000000000100000000000000010000000000000001000000000000,
        104'b00000000000000000000000000000000000100000000000000000000000000000000000000010000000000010000000000000000,
        104'b00000001000000000000000000000000000100000000000000000000001000000000000000000000000000010000000000000001,
        104'b00000000000000000000000000000000000100000001001000000000000000000000000000000000000000000000000000000000,
        104'b00000000000000000000000000100000000000000000001000000001000000000000000000000000000000000000000000000001,
        104'b00000000000000000000000000000001000100000000000100010000000100000000000000000000000000100000000000010010,
        104'b00000000000000010000000000000000000000000000000100010000000100010000000000000001000000100001000000000000,
        104'b00000000000000000000000000000000000100000000000100000000000000000000000000000000000000010001000000010000,
        104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010001,
        104'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000001,
        104'b00000000000000000000000000010000000000000001000000000000000000000000000000010000000000000000000000000001,
        104'b00000000000000000000000000000000000100000000000000010000000000000000000000000000000000000000000000000001,
        104'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000000000000000000000001000000000000000100000000000000010000000000010000000000000000,
        104'b00000000000000000000000100000001000100000000000100000000000000000000000000000000000000010000000100000000,
        104'b00000000000000000000000000010001000000000000000000010000000000010000000000010000000000000000000000000001,
        104'b00000000000000000000000100000001000000000000000000000000000000000000000000000000000000010000000000000000,
        104'b00000000000000000001000000000000000100000000000000000000000000000000000000000000000000010000000000010001,
        104'b00000000000000000000000100000000000000010000000000010000000000000000000000000000000000100000000000000000,
        104'b00000001000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000010000,
        104'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000100010000000000000000,
        104'b00000001000000000000000000010000000000000000000000000000000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000000000000000000000000000100010000000000000000000000000000000000000000000000000000,
        104'b00000001000000000000000100000001000000000000000000010000000000000000000000000000000000000001000000000001,
        104'b00000000000000000000000100000001000000000000000100000000000000000000000000010000000000010000000000000000,
        104'b00000001000000000000000100000000000000000000000000100000000000000000000000000000000100000000000000000000,
        104'b00000000000000000000000100000000000000000001000100000000000100000000000000000000000000010000000100000000,
        104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100100000000000010000,
        104'b00000000000000000000000000000001000100000010000000000000000000000000000000000000000000010000000000000010,
        104'b00000000000000000000000000000000001000000000000100010000000000000000000000000000000000010000000100000000,
        104'b00000001000000000000000000010000000000000000000000000000000000000000000000010000000000010000000000000000,
        104'b00000000000000000000000000010001000000000000000000000000000000000000000000010000000000100000000000000000,
        104'b00000000000000000000000000000001000000000000000100000000000000000000000000000000000000010001000000000000,
        104'b00000000000000010000000000000000000100000000000100000000000000000000000000000001000000000000000000000000,
        104'b00000000000000000000000000000001000000000001000000010000000000000000000000000000000000100010000000000000,
        104'b00000000000000000000000000000000000000000000000000000001000000010000000000000000000000010000000000000001,
        104'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000100001000000000000,
        104'b00000000000100000000000100010001000000000000000000000000000000000000000000010000000000100001000000000001,
        104'b00000000000000000000000000000001000000000000001000000000000100010000000000000000000000000000000000000000,
        104'b00000000000000000000000000000001000000000000000100010000000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000000010001000000000000000100000000000000000000000000010000000000000000000000000000,
        104'b00000000000000000000000100000000000100000000000100010000000000000000000000000000000000000001000000000001,
        104'b00000000000000000000000000000000000000000000000100000000000000000000000000000000001000100000000100000000,
        104'b00000000000000000001000000000000000000000000000000000000000000000000000000010000000000010000000000000001,
        104'b00000000000000000000000000010001000000000000000000000000000100000000000000000000000000000000000000000001,
        104'b00000000000000010000000000000000000000000000000100000000001000000000000000000000000000000000000000000001,
        104'b00000000000000000000000000000010000000000000000100000000000000000000000000000000000000000000000000010000,
        104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000000000000,
        104'b00000000000000000000000000010001000000000000000000000000000000010000000000000000000000010000000000000001,
        104'b00000000000000000000000000000001000000000000000000000000000100000000000000000000000100100000000000000000,
        104'b00000000000000010000000000000000000100000000000100010000000000000000000000000001000000000000000000000000,
        104'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000010000000000010000,
        104'b00000000000000000000000100010000000000000000000000000000000100000000000000000000000100000000000000000001,
        104'b00000000000000000000000100000000000100000000000100000000000000000000000000000000000000000000000000000000,
        104'b00000000000000000000000000010000000000000000000100000000000000000000000000000000000000000000000000000000,
        104'b00000000000000000000000100000000000100000000000000010000000000000000000000010000000000010010000000000000,
        104'b00000000000000000000000000000001000000000000001000000000000100000000000000010000000000000000000100000000,
        104'b00000000000000000000000100010000001000000000000000010000000000000000000000010010000000010010000000000010,
        104'b00000000000000000000000100010000000000000000000000000000000000000000000000000000000000010000000100000000,
        104'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100010001,
        104'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000001,
        104'b00000000000000000000000000000001000100000001000100010000000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000000000000000000000000000000010000000000010000000000000000000000010000000100000000,
        104'b00000001000000000000000000010000000100000000000100000000000000000000000000000000000100000000000000000000,
        104'b00000000000000000000000000000000000000000000001000000000000000010000000000000000000000000000000000010000,
        104'b00000000000000010000000000000001000000000000000000000000000100010000000000000000000000000000000000000001,
        104'b00000000000000000000000000000001000000000000001000000000000000000000000000000000000100010001000000000001,
        104'b00000001000000000000000000000000000000000000000000100000000000000000000000000000000000000000000100000001,
        104'b00000000000000000000000000000000000100000000000100000000000000000000000000010000000000010000000000000000,
        104'b00000001000000000000000000010000000100000001000000000000000000000000000000000000000000000000000000000001,
        104'b00000000000000000000000000010000001000000000000100010001000000000000000000010001000000010001000000000001,
        104'b00000001000000000000000000000000000100000000000000010000000000000000000000000001000000000000000000000001,
        104'b00000000000000000000000000000001000000000000000000000000000100000000000000000000000100010000000000000001,
        104'b00000000000000000000000000000000000100000000000100010000000000000000000000000000000000000000000000000000,
        104'b00000000000000010000000000000000000000000000000000010000000000000000000000010000000000010000000000000000,
        104'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000001,
        104'b00000000000000000000000000010000000000000000000000000000000100000000000000000000000000010000000000000001,
        104'b00000000000000000000000100000000000000000000000000010000000000000000000000000000000000000000000000010000,
        104'b00000000000000000000000000000000000000000000000100010001000100000000000000000000000000010000000000000000,
        104'b00000000000000000000000000000000001000000000000000010000000000000000000000000001000000010000000000000010,
        104'b00000000000000000000000000000000000100000000000000000000000000000000000000000001000000100000000000000001,
        104'b00000001000000000000000100000000001000000000000000000000000000000000000000010000000000000000000000000000,
        104'b00000000000000000000000000010000000000000000000000000000000000000000000000010000000000010001000000000001,
        104'b00000000000000000000000000010000000100000000000000000000000000000000000000010000000000100000000000000000,
        104'b00000000000000000000000100010000000100000000000100000000000100000000000000000000000000010000000000010000,
        104'b00000000000000000000000000000000000100000000000000010000000000000000000000000000000000010000000000000001,
        104'b00000000000000010000000100000000000000000000000100000000000100000000000000000000000000000001000000000000,
        104'b00000000000000000000000000100001000100000000000000000000000000000000000000000000000000000000000000000001,
        104'b00000000000000000000000100010001000000000000000000000000000000000000000000000001000000010000000000000000,
        104'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000010000000000000000,
        104'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000100000001000000000000,
        104'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000100000000000000000,
        104'b00000000000000000000000100100001000100000000000000000000000000000000000000000000000000000000000000000000,
        104'b00000000000000000000000000000001000000000000000000000001001000000000000000000000000000010000000000000000,
        104'b00000001000000000000000000000000000000000000000100010000000000000001000000000000000000010000000000000000,
        104'b00000000000000000001000000000000000100000000000100000000000000000000000000000000000100000000000000000001,
        104'b00000000000000000000000100000000000000000000000000000001000000000000000000000000000000000001000000010000,
        104'b00000000000000000000000000000001000100000000000000000000000000000000000000000000000000000001000100000001,
        104'b00000000000000000000000000000000000100000000000000000001000000000000000000000000000000010001000000000001,
        104'b00000000000000000000000000000000000000000000000100000000000100000000000000000000000000000000000100000001,
        104'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000001000000000001,
        104'b00000000000000010000000000000000000000000000000000010000000000000000000000000001000000000000000000000001,
        104'b00000000000000000000000000000000000000000010000000010000000000000000000000010000000000100001000000000001,
        104'b00000000000000010000000000000000000000000000000100010000000000010000000000000000000000000000000000000000,
        104'b00000000000000010000000000000000000000000000000000000000000100010000000000000000000000010001000000000001,
        104'b00000001000000000000000000000001000000000000000100010000000000000000000000000001000000010000000000010000,
        104'b00000000000000000000000000000001000000000000000000000000001000000000000000010000000000000000000000000001,
        104'b00000000000000000001000000000001000100000000000000000000000000000000000000000000000000100001000000000000,
        104'b00000000000000010000000000000000000000000000000000010000000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000100000001000000010000000000000000000100000000000000000000000000010000000000000001,
        104'b00000000000000000000000000010000000000000000000000000001000000000000000000000000000000010000000000000001,
        104'b00000000000000000000000000000000000000000010000000000000000100000000000000000000000000010000000000000001,
        104'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000010001000000000001,
        104'b00000000000000010000000000010000000000000000000000000000000000000000000000010000000000000000000000000001,
        104'b00000000000000000000000000010000000000000000000000000000000000010000000000000000000000010000000000000001,
        104'b00000000000000000000000000000000000000000000000100000000000100000000000000000000000000000001000100000000,
        104'b00000000000000000000000000000000000000000000000100000001000000000000000000010000000000010000000000000000,
        104'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000010000000000010000,
        104'b00000000000000000000000100000001000000000000000100010000000000000000000000000000000000000001000000000000,
        104'b00000000000000000000000000000000000000000000000000010001000000000000000000000000000000000000000000000001,
        104'b00000000000000000000000000010001000000000000000000010000000000000000000000000000000100010000000000000001,
        104'b00000000000000000000000000000000000000000001000000010000000100000000000000000000000000010000000000000001,
        104'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000010001000000000001,
        104'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001,
        104'b00000001000000000000000000000000000100000000000000000000000000000000000000000000000000010001000000000001,
        104'b00000000000000000000000000000010000000000000000000000001000000000000000000000000000000100000000000000000,
        104'b00000000000000000000000000010000000000000000000000010000000000000000000000010000000000000000000000000001,
        104'b00000000000000000000000100010000000000000000000100000000000000000000000000000000000000000000000000000000,
        104'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001,
        104'b00000001000000000000000000000001001000000000000100000000000000000000000000000000000000000000000000000000,
        104'b00000001000000000000000000000000000000000000000100010000000000000000000000000000000000010001000000010000,
        104'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000010001000000000010,
        104'b00000000000000000000000000000000000000000000000000000001000000000000000000010000000000000000000000000001,
        104'b00000000000000000000000000000000000000000000000000010000000000010000000000000000000000100000000000000000,
        104'b00000000000000000000000100000000000000000000000000010000000100000000000000000000000000010000000100000000,
        104'b00000000000000000000000000000000000100000001000100000001000100000000000000000000000000010000000000010000,
        104'b00000000000000000001000000000000000000000000000100000000000000000000000000000000000000010000000000010001,
        104'b00000000000000000000000000000000000000000000000000000001000100000000000000000000000000010000000000000001,
        104'b00000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000010,
        104'b00000001000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000001,
        104'b00000001000000000000000100000001000100000000000100000000000100000000000000000000000100010000000000000000,
        104'b00000000000000000000000000010000000000000001000000000000000000000000000000000000000000010000001000000001,
        104'b00000000000000010000000000010000000000000000000000000000000000000000000000010000000000000000000100000001,
        104'b00000000000000000000000100000000000000000000000100010000000000000000000000000000000100010010000000000000,
        104'b00000000000000010000000000000000000000000000000100010001000000000000000000000000000000000000000000000001,
        104'b00000000000000000000000000000000000000000001000000010000000000000001000000000000000000000000000000000010,
        104'b00000000000000000000000000000001000100000001000000000000000000000000000000010000000000000000000000000001,
        104'b00000000000000000000000000000000000000000000000100000000000000000000000000000000001000000000000000000000,
        104'b00000010000000000001000000000000000100000000000000000000000000000000000000000000000000100001000000000001,
        104'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000010001000100000001,
        104'b00000000000000000000000000000000000000000000000100100000000000000000000000000000000000010000000000000000,
        104'b00000001000000000000000000000000000000000001000000000000000100000000000000000000000000000000000000000001,
        104'b00000000000000000000000100010000000000000000000000000001000000000000000000010000000000000000000000010000,
        104'b00000000000000000000000000010000000000000000000000000000000100000000000000000000000000010000000000000000,
        104'b00000001000000000000000000000000000100000000000100000010000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000100000000000000000000,
        104'b00000000000000000000000000000000000000000000000100010000000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001000000000000,
        104'b00000000000000000000000100010000000100000000000000000000000000000000000000010001000000010001000000000001,
        104'b00000000000000000000000000010000000000000000000000000000001000000000000000000000000000010000000000000000,
        104'b00000000000000000000000000000000000000000000000100010000000100000000000000000001000000000000000000000000,
        104'b00000001000000000000000000000000000100000000000000000000000000000000000000000001000000100001000000000000,
        104'b00000000000000000000000000000000000100000000000100000000000000010000000000000000000000010000000000010000,
        104'b00000000000000000000000000100001000100000000000000000000000000000000000000000000000000100000000000000000,
        104'b00000000000000010000000000010000001000000000001100000001000000000000000000000000000000000000000000000000,
        104'b00000000000000000000000000000010000100000000000000000000000000000000000000000000000000100010000000000000,
        104'b00000000000000000000000000010000000000000000000000010000000000000000000000010000000000010000000000000000,
        104'b00000001000000010000000000000000001000000000000100000000000000000000000000000000000000000000000000000000,
        104'b00000000000000010000000000000000000000000000000100000000001000000000000000000000000100010000000000000000,
        104'b00000000000000000000000100000001000000000000000100000000000100000000000000000000000000000000000000000000,
        104'b00000000000000000000000000000000000000000000000100000000000100000000000000000001000000000000000000000001,
        104'b00000000000000000000000000000001000000000000000000000000000000000000000000010000000000110000000100000000,
        104'b00000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000001,
        104'b00000001000000000000000000000000001000000000000000000001000000000000000000000000000000000000000000000001,
        104'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000100000001,
        104'b00000000000000000000000000000000000100000000000100010000000000010000000000000000000000010000000000010000,
        104'b00000000000000000000000100000000000100000000000100000001000000000000000000010000000000000000000000000000,
        104'b00000000000000000000000000010000000000000000001000000000000000000000000000000000000100000000000000000000,
        104'b00000000000000010000000000000000000000000000000100000000000100000000000000000000000000010000000000010000,
        104'b00000000000000010000000000000010000100000000000000010000000000000000000000000000000000010000000000000001,
        104'b00000000000000000000000000000010000000000000000100010000000000000000000000000000000000010000000000000001,
        104'b00000000000000000000000100000000001000000000000100000001000000000000000000000000000000000000000000000000,
        104'b00000000000000000000000000010000000000000000000000010000000000000000000000000000000000010000000000000000,
        104'b00000000000000000000000000000001000000000000000100000000000000000000000000000000000000000000000000000000,
        104'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000001,
        104'b00000000000000000000000000000000000000000000000100010000000100000000000000000001000000000000000000000001,
        104'b00000000000000000000000100000001000000000000000100000001000000000000000000000000000100000000000000000001,
        104'b00000001000000000000000100000000000000000000000000000000000000000000000000000001000000000000000000000000,
        104'b00000000000000000000000000000000000000000000000100000000000000000001000000000000000000000000000000010000,
        104'b00000000000000000000000000010000001000000001000000010000000000000000000000000000000000010000000000000001,
        104'b00000000000000000000000000010000000100000000000000000000000000000000000000010000000100010000000000000001,
        104'b00000000000000000000000000000000000000000000001000000000000100010000000000000000000000000000000000000000,
        104'b00000000000000000000000000010001000000000000000000000000000000000000000000000000000000010000000000000001,
        104'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000100010000000000000000,
        104'b00000000000000000001000000000001000000000000000000010000000000000000000000000000000000100000000000000000,
        104'b00000000000000010000000000000000000000000000000000000000000000010000000000000000000000010000000000000001,
        104'b00000000000000000000000000000000000000000000000000000000000100000000000000010000000100000000000000000001,
        104'b00000001000000000000000000010000000000000000000100000000000000000000000000000000000000000001000000000001,
        104'b00000001000000000000000000000001000000000000000000000001000100000000000000000000000100010000000000000000,
        104'b00000000000000010000000000000000000000000000000000010000000000010000000000000000000000010000000000000000,
        104'b00000001000000000001000000000000000100000000000000000000000000000000000000000000000000100000000000000000,
        104'b00000000000000000000000000000000000100000000001000000000000100000000000000000000000000000000000100000000,
        104'b00000000000000000000000000000000000100000001000000000000000000000000000000000000000000010000000000000001,
        104'b00000001000000000000000100000001000100000000000100000000000000000000000000000000000000000000000000000000,
        104'b00000000000000000000000100000001000000000000000100000000000100000001000000000000000000010000000000000001,
        104'b00000000000000000000000000000001000000000000000100000001000000000000000000000000000000010000000000000000,
        104'b00000000000000010000000000000000000000000000001000000000001000000000000000000000000100000000000000000000,
        104'b00000000000000000000000100000000000100000000000100000000000100000000000000000000000100000000000000000000,
        104'b00000000000000000000001000100000000000000000000100000000000100000000000000100001000100000000000000000000,
        104'b00000000000000000000000000000000000000000000000000010001000000000000000000000000000000010000000000000001,
        104'b00000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000
	};
	
	localparam bit [7:0] alphabet [0:25] = '{
		8'b00000001,
		8'b00000010,
		8'b00000011,
		8'b00000100,
		8'b00000101,
		8'b00000110,
		8'b00000111,
		8'b00001000,
		8'b00001001,
		8'b00001010,
		8'b00001011,
		8'b00001100,
		8'b00001101,
		8'b00001110,
		8'b00001111,
		8'b00010000,
		8'b00010001,
		8'b00010010,
		8'b00010011,
		8'b00010100,
		8'b00010101,
		8'b00010110,
		8'b00010111,
		8'b00011000,
		8'b00011001,
		8'b00011010
	};
	
	// local parameters
	localparam S_IDLE      = 3'd0;
	localparam S_PRE_CALC  = 3'd1;
	localparam S_CALC      = 3'd2;
	localparam S_POST_CALC = 3'd3;
	localparam S_DONE      = 3'd4;
	
	// logics
	logic [2:0]              state_r, state_w;
	logic                    finish_r, finish_w;
	logic [COUNT_SIZE - 1:0] word_count_r, word_count_w;
	// logic [119:0]            word_r, word_w;
	// logic                    similarity_word_w  [0:COUNT_DICT_SIZE - 1], similarity_word_r  [0:COUNT_DICT_SIZE - 1];
    logic [9:0]              topN_similarity_w[0:19], topN_similarity_r[0:19];
    logic [14:0]             topN_value_w[0:19], topN_value_r[0:19];
    logic [9:0]              tmp_similarity_w[0:19], tmp_similarity_r[0:19];
    logic [14:0]             tmp_value_w[0:19], tmp_value_r[0:19];
	
	logic [3:0]              word_length_r, word_length_w;
    logic [3:0]              dict_word_length;
    logic [3:0]              prev_dict_word_length_r, prev_dict_word_length_w;
	
	logic [14:0]             similarity_value_w, similarity_value_r;
	logic [14:0]             max_similarity_value_r, max_similarity_value_w;
	logic [9:0]              wd_r, wd_w;
	logic [4:0]              ptr_r, ptr_w;
	
	// integer i, j, ptr_word;
	
	// assign values
	assign o_similarity_finish = finish_r;
	assign o_similarity_word = topN_similarity_r;
    assign dict_word_length = count_dict[wd_r][3:0] + count_dict[wd_r][7:4] + count_dict[wd_r][11:8] + count_dict[wd_r][15:12] + count_dict[wd_r][19:16] + count_dict[wd_r][23:20] + count_dict[wd_r][27:24] + count_dict[wd_r][31:28] + count_dict[wd_r][35:32] + count_dict[wd_r][39:36] + count_dict[wd_r][43:40] + count_dict[wd_r][47:44] + count_dict[wd_r][51:48] + count_dict[wd_r][55:52] + count_dict[wd_r][59:56] + count_dict[wd_r][63:60] + count_dict[wd_r][67:64] + count_dict[wd_r][71:68] + count_dict[wd_r][75:72] + count_dict[wd_r][79:76] + count_dict[wd_r][83:80] + count_dict[wd_r][87:84] + count_dict[wd_r][91:88] + count_dict[wd_r][95:92] + count_dict[wd_r][99:96] + count_dict[wd_r][103:100];

	always_comb begin
		state_w = state_r;
		finish_w = finish_r;
		word_count_w = word_count_r;
		// word_w = word_r;
		similarity_value_w = similarity_value_r;
		max_similarity_value_w = max_similarity_value_r;
		wd_w = wd_r;
		ptr_w = ptr_r;
		word_length_w = word_length_r;

        prev_dict_word_length_w = prev_dict_word_length_r;

        topN_similarity_w = topN_similarity_r;
        topN_value_w = topN_value_r;
        tmp_similarity_w = tmp_similarity_r;
        tmp_value_w = tmp_value_r;
		
		case (state_r)
			S_IDLE: begin
				finish_w = 1'b0;
				if (i_similarity_start) begin
					state_w = S_PRE_CALC;
                    similarity_value_w = 0;
                    topN_similarity_w = '{20{10'b0}};
                    topN_value_w = '{20{15'b0}};
                    tmp_similarity_w = '{20{10'b0}};
                    tmp_value_w = '{20{15'b0}};
				end
			end
			S_PRE_CALC: begin
				// calculate word length
                word_length_w = (i_similarity_word[7:0] != 8'b0) + (i_similarity_word[15:8] != 8'b0) + (i_similarity_word[23:16] != 8'b0) + (i_similarity_word[31:24] != 8'b0) + (i_similarity_word[39:32] != 8'b0) + (i_similarity_word[47:40] != 8'b0) + (i_similarity_word[55:48] != 8'b0) + (i_similarity_word[63:56] != 8'b0) + (i_similarity_word[71:64] != 8'b0) + (i_similarity_word[79:72] != 8'b0) + (i_similarity_word[87:80] != 8'b0) + (i_similarity_word[95:88] != 8'b0) + (i_similarity_word[103:96] != 8'b0) + (i_similarity_word[111:104] != 8'b0) + (i_similarity_word[119:112] != 8'b0);
				// $display(word_length_w);
				// $display(dict_word_length_w[399]);
                word_count_w = ((1 << ((i_similarity_word[4:0]) * 4)) + (1 << ((i_similarity_word[12:8]) * 4)) + (1 << ((i_similarity_word[20:16]) * 4)) + (1 << ((i_similarity_word[28:24]) * 4)) + (1 << ((i_similarity_word[36:32]) * 4)) + (1 << ((i_similarity_word[44:40]) * 4)) + (1 << ((i_similarity_word[52:48]) * 4)) + (1 << ((i_similarity_word[60:56]) * 4)) + (1 << ((i_similarity_word[68:64]) * 4)) + (1 << ((i_similarity_word[76:72]) * 4)) + (1 << ((i_similarity_word[84:80]) * 4)) + (1 << ((i_similarity_word[92:88]) * 4)) + (1 << ((i_similarity_word[100:96]) * 4)) + (1 << ((i_similarity_word[108:104]) * 4)) + (1 << ((i_similarity_word[116:112]) * 4))) >> 4;
                // similarity_value_w = (word_count_r[3:0] * count_dict[wd_r][3:0]) + (word_count_r[7:4] * count_dict[wd_r][7:4]) + (word_count_r[11:8] * count_dict[wd_r][11:8]) + (word_count_r[15:12] * count_dict[wd_r][15:12]) + (word_count_r[19:16] * count_dict[wd_r][19:16]) + (word_count_r[23:20] * count_dict[wd_r][23:20]) + (word_count_r[27:24] * count_dict[wd_r][27:24]) + (word_count_r[31:28] * count_dict[wd_r][31:28]) + (word_count_r[35:32] * count_dict[wd_r][35:32]) + (word_count_r[39:36] * count_dict[wd_r][39:36]) + (word_count_r[43:40] * count_dict[wd_r][43:40]) + (word_count_r[47:44] * count_dict[wd_r][47:44]) + (word_count_r[51:48] * count_dict[wd_r][51:48]) + (word_count_r[55:52] * count_dict[wd_r][55:52]) + (word_count_r[59:56] * count_dict[wd_r][59:56]) + (word_count_r[63:60] * count_dict[wd_r][63:60]) + (word_count_r[67:64] * count_dict[wd_r][67:64]) + (word_count_r[71:68] * count_dict[wd_r][71:68]) + (word_count_r[75:72] * count_dict[wd_r][75:72]) + (word_count_r[79:76] * count_dict[wd_r][79:76]) + (word_count_r[83:80] * count_dict[wd_r][83:80]) + (word_count_r[87:84] * count_dict[wd_r][87:84]) + (word_count_r[91:88] * count_dict[wd_r][91:88]) + (word_count_r[95:92] * count_dict[wd_r][95:92]) + (word_count_r[99:96] * count_dict[wd_r][99:96]) + (word_count_r[103:100] * count_dict[wd_r][103:100]);
				// tmp_similarity_w[0] = 0;
                wd_w = 0;
				state_w = S_CALC;
			end
			S_CALC: begin
				// calculate each similarity value
				if (wd_r == COUNT_DICT_SIZE - 1 + 20) begin
					state_w = S_DONE;
				end else begin
                    if (wd_r < COUNT_DICT_SIZE) begin
                        similarity_value_w = (word_count_r[3:0] * count_dict[wd_r][3:0]) + (word_count_r[7:4] * count_dict[wd_r][7:4]) + (word_count_r[11:8] * count_dict[wd_r][11:8]) + (word_count_r[15:12] * count_dict[wd_r][15:12]) + (word_count_r[19:16] * count_dict[wd_r][19:16]) + (word_count_r[23:20] * count_dict[wd_r][23:20]) + (word_count_r[27:24] * count_dict[wd_r][27:24]) + (word_count_r[31:28] * count_dict[wd_r][31:28]) + (word_count_r[35:32] * count_dict[wd_r][35:32]) + (word_count_r[39:36] * count_dict[wd_r][39:36]) + (word_count_r[43:40] * count_dict[wd_r][43:40]) + (word_count_r[47:44] * count_dict[wd_r][47:44]) + (word_count_r[51:48] * count_dict[wd_r][51:48]) + (word_count_r[55:52] * count_dict[wd_r][55:52]) + (word_count_r[59:56] * count_dict[wd_r][59:56]) + (word_count_r[63:60] * count_dict[wd_r][63:60]) + (word_count_r[67:64] * count_dict[wd_r][67:64]) + (word_count_r[71:68] * count_dict[wd_r][71:68]) + (word_count_r[75:72] * count_dict[wd_r][75:72]) + (word_count_r[79:76] * count_dict[wd_r][79:76]) + (word_count_r[83:80] * count_dict[wd_r][83:80]) + (word_count_r[87:84] * count_dict[wd_r][87:84]) + (word_count_r[91:88] * count_dict[wd_r][91:88]) + (word_count_r[95:92] * count_dict[wd_r][95:92]) + (word_count_r[99:96] * count_dict[wd_r][99:96]) + (word_count_r[103:100] * count_dict[wd_r][103:100]);
                        tmp_similarity_w[0] = wd_r - 1;
                        prev_dict_word_length_w = dict_word_length;
                        if (word_length_r <= prev_dict_word_length_r) begin
                            tmp_value_w[0] = (similarity_value_r << 10) / prev_dict_word_length_r;
                        end else begin
                            tmp_value_w[0] = (similarity_value_r << 10) / word_length_r;
                        end
                    end
                    else begin
                        tmp_value_w[0] = 0;
                    end

                    // $display("%d, %d", wd_r - 1, similarity_value_r);

                    for (integer i = 0; i < 19; i = i + 1) begin
                        if (tmp_value_r[i] > topN_value_r[i]) begin
                            topN_value_w[i] = tmp_value_r[i];
                            topN_similarity_w[i] = tmp_similarity_r[i];
                            tmp_value_w[i+1] = topN_value_r[i];
                            tmp_similarity_w[i+1] = topN_similarity_r[i];
                        end else begin
                            tmp_value_w[i+1] = tmp_value_r[i];
                            tmp_similarity_w[i+1] = tmp_similarity_r[i];
                        end
                    end

                    if (tmp_value_r[19] > topN_value_r[19]) begin
                        topN_value_w[19] = tmp_value_r[19];
                        topN_similarity_w[19] = tmp_similarity_r[19];
                    end
					

					// if (similarity_value_w[wd_r] >= max_similarity_value_r) begin
					// 	max_similarity_value_w = similarity_value_w[wd_r];
					// end
					wd_w = wd_r + 1;
				end
			end
			// S_POST_CALC: begin
			// 	// find the biggest 20 values
			// 	if (ptr_r >= 20) begin
			// 		state_w = S_DONE;
			// 	end else begin
			// 		for (ptr_word = 0; ptr_word < COUNT_DICT_SIZE; ptr_word = ptr_word + 1) begin
			// 			if (ptr_w >= 20) begin
			// 				break;
			// 			end
			// 			if (similarity_value_w[ptr_word] == max_similarity_value_r) begin
			// 				similarity_word_w[ptr_word] = 1'b1;
			// 				ptr_w = ptr_w + 1;
			// 			end
			// 		end
			// 	end
				
			// 	max_similarity_value_w = max_similarity_value_r - 5'd1;
			// end
			S_DONE: begin
				finish_w = 1'b1;
				state_w = S_IDLE;
			end
		endcase
		
	end

	always_ff @ (posedge i_similarity_clk or posedge i_similarity_rst_n) begin
		if (i_similarity_rst_n) begin
			state_r                <= S_IDLE;
			finish_r               <= 1'b0;
			word_count_r           <= 104'b0;
			// word_r                 <= 120'b0;
			// similarity_word_r      <= '{500{1'b0}};
			similarity_value_r     <= 15'b0;
			max_similarity_value_r <= 15'b0;
			wd_r                   <= 9'b0;
			ptr_r                  <= 5'b0;
			word_length_r          <= 4'b0;
            prev_dict_word_length_r <= 4'b0;
			// dict_word_length_r     <= '{500{4'b0}};

            topN_similarity_r <= '{20{10'b0}};
            topN_value_r <= '{20{15'b0}};
            tmp_similarity_r <= '{20{10'b0}};
            tmp_value_r <= '{20{15'b0}};

		end else begin
			state_r                <= state_w;
			finish_r               <= finish_w;
			word_count_r           <= word_count_w;
			// word_r                 <= word_w;
			// similarity_word_r      <= similarity_word_w;
			similarity_value_r     <= similarity_value_w;
			max_similarity_value_r <= max_similarity_value_w;
			wd_r                   <= wd_w;
			ptr_r                  <= ptr_w;
			word_length_r          <= word_length_w;
            prev_dict_word_length_r <= prev_dict_word_length_w;
			// dict_word_length_r     <= dict_word_length_w;

            topN_similarity_r <= topN_similarity_w;
            topN_value_r <= topN_value_w;
            tmp_similarity_r <= tmp_similarity_w;
            tmp_value_r <= tmp_value_w;
		end
	end
endmodule

`timescale 1ns / 100ps

module tb;
    localparam CLK = 10;
    localparam HCLK = CLK / 2;
    localparam SF = 2.0 ** -8.0;

    localparam bit [119:0] DTW_candidate_word [0:19] = '{
        120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000100110001000000011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000100100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000111100000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110001000000000111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101000000100000100100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001101000000011,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100000010100000100100010101,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001000101010000101000011000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100001000000011010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100001010,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010001000000001111,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100010000,
		120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000011
    };

    logic clk, rst, start, finished, valid;
    logic [2:0] state;
    logic [4:0] word_num;
    logic [14:0] dp;
    logic [119:0] word_in = 120'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100010001;
    logic [119:0] word_out;

    initial clk = 0;
    always #HCLK clk = ~clk;

    DTW dtw1 (
        .i_DTW_clk(clk),
        .i_DTW_rst_n(rst),
        .i_DTW_start(start),
        .i_DTW_word(word_in),
        .i_DTW_candidate_word(DTW_candidate_word),
        .o_DTW_finish(finished),
        .o_DTW_word(word_out),
        .o_state(state)
    );

    initial begin
        $fsdbDumpfile("final.fsdb");
        $fsdbDumpvars;

        rst <= 0;
        start <= 0;
        #(2 * CLK);
        rst <= 1;
        @(posedge clk) rst <= 0;

        $display("==========input=============");
        $display("%b", word_in);

        start <= 1;
        #(CLK)
        start <= 0;
        // #(10 * CLK);

        while (!finished) begin
            // $display(word_length);
            #(CLK);
        end
        $display();
        $display("==========output=============");
        $display("%b", word_out);
        $finish;
    end

    initial begin
		#(5000000*CLK)
		$display("Too Slow, Abort");
		$finish;
	end

endmodule